--------------------------------------------------------------------------------
-- Company: <Name>
--
-- File: Index_rom.vhd
-- File history:
--      <Revision number>: <Date>: <Comments>
--      <Revision number>: <Date>: <Comments>
--      <Revision number>: <Date>: <Comments>
--
-- Description: 
--
-- <Description here>
--
-- Targeted device: <Family::PolarFire> <Die::MPF300T> <Package::FCG484>
-- Author: <Name>
--
--------------------------------------------------------------------------------

library IEEE;

use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;  -- 添加数值转换库
use IEEE.STD_LOGIC_UNSIGNED.ALL;
entity Index_rom is
port (
	clk : IN  std_logic; -- example
	rstn: IN  std_logic;
    address_in1 : in std_logic_vector(15 downto 0)  ;
	address_out1: out std_logic_vector(15 downto 0)  ;
	address_out2 : out std_logic_vector(15 downto 0) 
);
end Index_rom;
architecture architecture_Index_rom of Index_rom is
	type data_array is array(8919 downto 0)of std_logic_vector(15 downto 0);	
	constant rom_reg:data_array:=		
		(X"0004",
		X"00AB",
		X"012C",
		X"01D3",
		X"0254",
		X"02FB",
		X"037C",
		X"0423",
		X"04A4",
		X"054B",
		X"05CC",
		X"0673",
		X"06F4",
		X"079B",
		X"081C",
		X"08C3",
		X"0944",
		X"09EB",
		X"0A6C",
		X"0B13",
		X"0B94",
		X"0C3B",
		X"0CBC",
		X"0D63",
		X"0DE4",
		X"0E8B",
		X"0F0C",
		X"0FB3",
		X"1034",
		X"10DB",
		X"115C",
		X"1203",
		X"1284",
		X"132B",
		X"13AC",
		X"1453",
		X"14D4",
		X"157B",
		X"15FC",
		X"16A3",
		X"1724",
		X"17CB",
		X"184C",
		X"18F3",
		X"1974",
		X"1A1B",
		X"1A9C",
		X"1B43",
		X"1BC4",
		X"1C6B",
		X"1CEC",
		X"1D93",
		X"1E14",
		X"1EBB",
		X"1F3C",
		X"1FE3",
		X"2064",
		X"210B",
		X"218C",
		X"2233",
		X"22B4",
		X"0083",
		X"0104",
		X"01AB",
		X"022C",
		X"02D3",
		X"0354",
		X"03FB",
		X"047C",
		X"0523",
		X"05A4",
		X"064B",
		X"06CC",
		X"0773",
		X"07F4",
		X"089B",
		X"091C",
		X"09C3",
		X"0A44",
		X"0AEB",
		X"0B6C",
		X"0C13",
		X"0C94",
		X"0D3B",
		X"0DBC",
		X"0E63",
		X"0EE4",
		X"0F8B",
		X"100C",
		X"10B3",
		X"1134",
		X"11DB",
		X"125C",
		X"1303",
		X"1384",
		X"142B",
		X"14AC",
		X"1553",
		X"15D4",
		X"167B",
		X"16FC",
		X"17A3",
		X"1824",
		X"18CB",
		X"194C",
		X"19F3",
		X"1A74",
		X"1B1B",
		X"1B9C",
		X"1C43",
		X"1CC4",
		X"1D6B",
		X"1DEC",
		X"1E93",
		X"1F14",
		X"1FBB",
		X"203C",
		X"20E3",
		X"2164",
		X"220B",
		X"228C",
		X"005B",
		X"00DC",
		X"0183",
		X"0204",
		X"02AB",
		X"032C",
		X"03D3",
		X"0454",
		X"04FB",
		X"057C",
		X"0623",
		X"06A4",
		X"074B",
		X"07CC",
		X"0873",
		X"08F4",
		X"099B",
		X"0A1C",
		X"0AC3",
		X"0B44",
		X"0BEB",
		X"0C6C",
		X"0D13",
		X"0D94",
		X"0E3B",
		X"0EBC",
		X"0F63",
		X"0FE4",
		X"108B",
		X"110C",
		X"11B3",
		X"1234",
		X"12DB",
		X"135C",
		X"1403",
		X"1484",
		X"152B",
		X"15AC",
		X"1653",
		X"16D4",
		X"177B",
		X"17FC",
		X"18A3",
		X"1924",
		X"19CB",
		X"1A4C",
		X"1AF3",
		X"1B74",
		X"1C1B",
		X"1C9C",
		X"1D43",
		X"1DC4",
		X"1E6B",
		X"1EEC",
		X"1F93",
		X"2014",
		X"20BB",
		X"213C",
		X"21E3",
		X"2264",
		X"0033",
		X"00B4",
		X"015B",
		X"01DC",
		X"0283",
		X"0304",
		X"03AB",
		X"042C",
		X"04D3",
		X"0554",
		X"05FB",
		X"067C",
		X"0723",
		X"07A4",
		X"084B",
		X"08CC",
		X"0973",
		X"09F4",
		X"0A9B",
		X"0B1C",
		X"0BC3",
		X"0C44",
		X"0CEB",
		X"0D6C",
		X"0E13",
		X"0E94",
		X"0F3B",
		X"0FBC",
		X"1063",
		X"10E4",
		X"118B",
		X"120C",
		X"12B3",
		X"1334",
		X"13DB",
		X"145C",
		X"1503",
		X"1584",
		X"162B",
		X"16AC",
		X"1753",
		X"17D4",
		X"187B",
		X"18FC",
		X"19A3",
		X"1A24",
		X"1ACB",
		X"1B4C",
		X"1BF3",
		X"1C74",
		X"1D1B",
		X"1D9C",
		X"1E43",
		X"1EC4",
		X"1F6B",
		X"1FEC",
		X"2093",
		X"2114",
		X"21BB",
		X"223C",
		X"000B",
		X"008C",
		X"0133",
		X"01B4",
		X"025B",
		X"02DC",
		X"0383",
		X"0404",
		X"04AB",
		X"052C",
		X"05D3",
		X"0654",
		X"06FB",
		X"077C",
		X"0823",
		X"08A4",
		X"094B",
		X"09CC",
		X"0A73",
		X"0AF4",
		X"0B9B",
		X"0C1C",
		X"0CC3",
		X"0D44",
		X"0DEB",
		X"0E6C",
		X"0F13",
		X"0F94",
		X"103B",
		X"10BC",
		X"1163",
		X"11E4",
		X"128B",
		X"130C",
		X"13B3",
		X"1434",
		X"14DB",
		X"155C",
		X"1603",
		X"1684",
		X"172B",
		X"17AC",
		X"1853",
		X"18D4",
		X"197B",
		X"19FC",
		X"1AA3",
		X"1B24",
		X"1BCB",
		X"1C4C",
		X"1CF3",
		X"1D74",
		X"1E1B",
		X"1E9C",
		X"1F43",
		X"1FC4",
		X"206B",
		X"20EC",
		X"2193",
		X"2214",
		X"22BB",
		X"0064",
		X"010B",
		X"018C",
		X"0233",
		X"02B4",
		X"035B",
		X"03DC",
		X"0483",
		X"0504",
		X"05AB",
		X"062C",
		X"06D3",
		X"0754",
		X"07FB",
		X"087C",
		X"0923",
		X"09A4",
		X"0A4B",
		X"0ACC",
		X"0B73",
		X"0BF4",
		X"0C9B",
		X"0D1C",
		X"0DC3",
		X"0E44",
		X"0EEB",
		X"0F6C",
		X"1013",
		X"1094",
		X"113B",
		X"11BC",
		X"1263",
		X"12E4",
		X"138B",
		X"140C",
		X"14B3",
		X"1534",
		X"15DB",
		X"165C",
		X"1703",
		X"1784",
		X"182B",
		X"18AC",
		X"1953",
		X"19D4",
		X"1A7B",
		X"1AFC",
		X"1BA3",
		X"1C24",
		X"1CCB",
		X"1D4C",
		X"1DF3",
		X"1E74",
		X"1F1B",
		X"1F9C",
		X"2043",
		X"20C4",
		X"216B",
		X"21EC",
		X"2293",
		X"003C",
		X"00E3",
		X"0164",
		X"020B",
		X"028C",
		X"0333",
		X"03B4",
		X"045B",
		X"04DC",
		X"0583",
		X"0604",
		X"06AB",
		X"072C",
		X"07D3",
		X"0854",
		X"08FB",
		X"097C",
		X"0A23",
		X"0AA4",
		X"0B4B",
		X"0BCC",
		X"0C73",
		X"0CF4",
		X"0D9B",
		X"0E1C",
		X"0EC3",
		X"0F44",
		X"0FEB",
		X"106C",
		X"1113",
		X"1194",
		X"123B",
		X"12BC",
		X"1363",
		X"13E4",
		X"148B",
		X"150C",
		X"15B3",
		X"1634",
		X"16DB",
		X"175C",
		X"1803",
		X"1884",
		X"192B",
		X"19AC",
		X"1A53",
		X"1AD4",
		X"1B7B",
		X"1BFC",
		X"1CA3",
		X"1D24",
		X"1DCB",
		X"1E4C",
		X"1EF3",
		X"1F74",
		X"201B",
		X"209C",
		X"2143",
		X"21C4",
		X"226B",
		X"0014",
		X"00BB",
		X"013C",
		X"01E3",
		X"0264",
		X"030B",
		X"038C",
		X"0433",
		X"04B4",
		X"055B",
		X"05DC",
		X"0683",
		X"0704",
		X"07AB",
		X"082C",
		X"08D3",
		X"0954",
		X"09FB",
		X"0A7C",
		X"0B23",
		X"0BA4",
		X"0C4B",
		X"0CCC",
		X"0D73",
		X"0DF4",
		X"0E9B",
		X"0F1C",
		X"0FC3",
		X"1044",
		X"10EB",
		X"116C",
		X"1213",
		X"1294",
		X"133B",
		X"13BC",
		X"1463",
		X"14E4",
		X"158B",
		X"160C",
		X"16B3",
		X"1734",
		X"17DB",
		X"185C",
		X"1903",
		X"1984",
		X"1A2B",
		X"1AAC",
		X"1B53",
		X"1BD4",
		X"1C7B",
		X"1CFC",
		X"1DA3",
		X"1E24",
		X"1ECB",
		X"1F4C",
		X"1FF3",
		X"2074",
		X"211B",
		X"219C",
		X"2243",
		X"22C4",
		X"0093",
		X"0114",
		X"01BB",
		X"023C",
		X"02E3",
		X"0364",
		X"040B",
		X"048C",
		X"0533",
		X"05B4",
		X"065B",
		X"06DC",
		X"0783",
		X"0804",
		X"08AB",
		X"092C",
		X"09D3",
		X"0A54",
		X"0AFB",
		X"0B7C",
		X"0C23",
		X"0CA4",
		X"0D4B",
		X"0DCC",
		X"0E73",
		X"0EF4",
		X"0F9B",
		X"101C",
		X"10C3",
		X"1144",
		X"11EB",
		X"126C",
		X"1313",
		X"1394",
		X"143B",
		X"14BC",
		X"1563",
		X"15E4",
		X"168B",
		X"170C",
		X"17B3",
		X"1834",
		X"18DB",
		X"195C",
		X"1A03",
		X"1A84",
		X"1B2B",
		X"1BAC",
		X"1C53",
		X"1CD4",
		X"1D7B",
		X"1DFC",
		X"1EA3",
		X"1F24",
		X"1FCB",
		X"204C",
		X"20F3",
		X"2174",
		X"221B",
		X"229C",
		X"006B",
		X"00EC",
		X"0193",
		X"0214",
		X"02BB",
		X"033C",
		X"03E3",
		X"0464",
		X"050B",
		X"058C",
		X"0633",
		X"06B4",
		X"075B",
		X"07DC",
		X"0883",
		X"0904",
		X"09AB",
		X"0A2C",
		X"0AD3",
		X"0B54",
		X"0BFB",
		X"0C7C",
		X"0D23",
		X"0DA4",
		X"0E4B",
		X"0ECC",
		X"0F73",
		X"0FF4",
		X"109B",
		X"111C",
		X"11C3",
		X"1244",
		X"12EB",
		X"136C",
		X"1413",
		X"1494",
		X"153B",
		X"15BC",
		X"1663",
		X"16E4",
		X"178B",
		X"180C",
		X"18B3",
		X"1934",
		X"19DB",
		X"1A5C",
		X"1B03",
		X"1B84",
		X"1C2B",
		X"1CAC",
		X"1D53",
		X"1DD4",
		X"1E7B",
		X"1EFC",
		X"1FA3",
		X"2024",
		X"20CB",
		X"214C",
		X"21F3",
		X"2274",
		X"0043",
		X"00C4",
		X"016B",
		X"01EC",
		X"0293",
		X"0314",
		X"03BB",
		X"043C",
		X"04E3",
		X"0564",
		X"060B",
		X"068C",
		X"0733",
		X"07B4",
		X"085B",
		X"08DC",
		X"0983",
		X"0A04",
		X"0AAB",
		X"0B2C",
		X"0BD3",
		X"0C54",
		X"0CFB",
		X"0D7C",
		X"0E23",
		X"0EA4",
		X"0F4B",
		X"0FCC",
		X"1073",
		X"10F4",
		X"119B",
		X"121C",
		X"12C3",
		X"1344",
		X"13EB",
		X"146C",
		X"1513",
		X"1594",
		X"163B",
		X"16BC",
		X"1763",
		X"17E4",
		X"188B",
		X"190C",
		X"19B3",
		X"1A34",
		X"1ADB",
		X"1B5C",
		X"1C03",
		X"1C84",
		X"1D2B",
		X"1DAC",
		X"1E53",
		X"1ED4",
		X"1F7B",
		X"1FFC",
		X"20A3",
		X"2124",
		X"21CB",
		X"224C",
		X"001B",
		X"009C",
		X"0143",
		X"01C4",
		X"026B",
		X"02EC",
		X"0393",
		X"0414",
		X"04BB",
		X"053C",
		X"05E3",
		X"0664",
		X"070B",
		X"078C",
		X"0833",
		X"08B4",
		X"095B",
		X"09DC",
		X"0A83",
		X"0B04",
		X"0BAB",
		X"0C2C",
		X"0CD3",
		X"0D54",
		X"0DFB",
		X"0E7C",
		X"0F23",
		X"0FA4",
		X"104B",
		X"10CC",
		X"1173",
		X"11F4",
		X"129B",
		X"131C",
		X"13C3",
		X"1444",
		X"14EB",
		X"156C",
		X"1613",
		X"1694",
		X"173B",
		X"17BC",
		X"1863",
		X"18E4",
		X"198B",
		X"1A0C",
		X"1AB3",
		X"1B34",
		X"1BDB",
		X"1C5C",
		X"1D03",
		X"1D84",
		X"1E2B",
		X"1EAC",
		X"1F53",
		X"1FD4",
		X"207B",
		X"20FC",
		X"21A3",
		X"2224",
		X"22CB",
		X"0074",
		X"011B",
		X"019C",
		X"0243",
		X"02C4",
		X"036B",
		X"03EC",
		X"0493",
		X"0514",
		X"05BB",
		X"063C",
		X"06E3",
		X"0764",
		X"080B",
		X"088C",
		X"0933",
		X"09B4",
		X"0A5B",
		X"0ADC",
		X"0B83",
		X"0C04",
		X"0CAB",
		X"0D2C",
		X"0DD3",
		X"0E54",
		X"0EFB",
		X"0F7C",
		X"1023",
		X"10A4",
		X"114B",
		X"11CC",
		X"1273",
		X"12F4",
		X"139B",
		X"141C",
		X"14C3",
		X"1544",
		X"15EB",
		X"166C",
		X"1713",
		X"1794",
		X"183B",
		X"18BC",
		X"1963",
		X"19E4",
		X"1A8B",
		X"1B0C",
		X"1BB3",
		X"1C34",
		X"1CDB",
		X"1D5C",
		X"1E03",
		X"1E84",
		X"1F2B",
		X"1FAC",
		X"2053",
		X"20D4",
		X"217B",
		X"21FC",
		X"22A3",
		X"004C",
		X"00F3",
		X"0174",
		X"021B",
		X"029C",
		X"0343",
		X"03C4",
		X"046B",
		X"04EC",
		X"0593",
		X"0614",
		X"06BB",
		X"073C",
		X"07E3",
		X"0864",
		X"090B",
		X"098C",
		X"0A33",
		X"0AB4",
		X"0B5B",
		X"0BDC",
		X"0C83",
		X"0D04",
		X"0DAB",
		X"0E2C",
		X"0ED3",
		X"0F54",
		X"0FFB",
		X"107C",
		X"1123",
		X"11A4",
		X"124B",
		X"12CC",
		X"1373",
		X"13F4",
		X"149B",
		X"151C",
		X"15C3",
		X"1644",
		X"16EB",
		X"176C",
		X"1813",
		X"1894",
		X"193B",
		X"19BC",
		X"1A63",
		X"1AE4",
		X"1B8B",
		X"1C0C",
		X"1CB3",
		X"1D34",
		X"1DDB",
		X"1E5C",
		X"1F03",
		X"1F84",
		X"202B",
		X"20AC",
		X"2153",
		X"21D4",
		X"227B",
		X"0024",
		X"00CB",
		X"014C",
		X"01F3",
		X"0274",
		X"031B",
		X"039C",
		X"0443",
		X"04C4",
		X"056B",
		X"05EC",
		X"0693",
		X"0714",
		X"07BB",
		X"083C",
		X"08E3",
		X"0964",
		X"0A0B",
		X"0A8C",
		X"0B33",
		X"0BB4",
		X"0C5B",
		X"0CDC",
		X"0D83",
		X"0E04",
		X"0EAB",
		X"0F2C",
		X"0FD3",
		X"1054",
		X"10FB",
		X"117C",
		X"1223",
		X"12A4",
		X"134B",
		X"13CC",
		X"1473",
		X"14F4",
		X"159B",
		X"161C",
		X"16C3",
		X"1744",
		X"17EB",
		X"186C",
		X"1913",
		X"1994",
		X"1A3B",
		X"1ABC",
		X"1B63",
		X"1BE4",
		X"1C8B",
		X"1D0C",
		X"1DB3",
		X"1E34",
		X"1EDB",
		X"1F5C",
		X"2003",
		X"2084",
		X"212B",
		X"21AC",
		X"2253",
		X"22D4",
		X"00A3",
		X"0124",
		X"01CB",
		X"024C",
		X"02F3",
		X"0374",
		X"041B",
		X"049C",
		X"0543",
		X"05C4",
		X"066B",
		X"06EC",
		X"0793",
		X"0814",
		X"08BB",
		X"093C",
		X"09E3",
		X"0A64",
		X"0B0B",
		X"0B8C",
		X"0C33",
		X"0CB4",
		X"0D5B",
		X"0DDC",
		X"0E83",
		X"0F04",
		X"0FAB",
		X"102C",
		X"10D3",
		X"1154",
		X"11FB",
		X"127C",
		X"1323",
		X"13A4",
		X"144B",
		X"14CC",
		X"1573",
		X"15F4",
		X"169B",
		X"171C",
		X"17C3",
		X"1844",
		X"18EB",
		X"196C",
		X"1A13",
		X"1A94",
		X"1B3B",
		X"1BBC",
		X"1C63",
		X"1CE4",
		X"1D8B",
		X"1E0C",
		X"1EB3",
		X"1F34",
		X"1FDB",
		X"205C",
		X"2103",
		X"2184",
		X"222B",
		X"22AC",
		X"007B",
		X"00FC",
		X"01A3",
		X"0224",
		X"02CB",
		X"034C",
		X"03F3",
		X"0474",
		X"051B",
		X"059C",
		X"0643",
		X"06C4",
		X"076B",
		X"07EC",
		X"0893",
		X"0914",
		X"09BB",
		X"0A3C",
		X"0AE3",
		X"0B64",
		X"0C0B",
		X"0C8C",
		X"0D33",
		X"0DB4",
		X"0E5B",
		X"0EDC",
		X"0F83",
		X"1004",
		X"10AB",
		X"112C",
		X"11D3",
		X"1254",
		X"12FB",
		X"137C",
		X"1423",
		X"14A4",
		X"154B",
		X"15CC",
		X"1673",
		X"16F4",
		X"179B",
		X"181C",
		X"18C3",
		X"1944",
		X"19EB",
		X"1A6C",
		X"1B13",
		X"1B94",
		X"1C3B",
		X"1CBC",
		X"1D63",
		X"1DE4",
		X"1E8B",
		X"1F0C",
		X"1FB3",
		X"2034",
		X"20DB",
		X"215C",
		X"2203",
		X"2284",
		X"0053",
		X"00D4",
		X"017B",
		X"01FC",
		X"02A3",
		X"0324",
		X"03CB",
		X"044C",
		X"04F3",
		X"0574",
		X"061B",
		X"069C",
		X"0743",
		X"07C4",
		X"086B",
		X"08EC",
		X"0993",
		X"0A14",
		X"0ABB",
		X"0B3C",
		X"0BE3",
		X"0C64",
		X"0D0B",
		X"0D8C",
		X"0E33",
		X"0EB4",
		X"0F5B",
		X"0FDC",
		X"1083",
		X"1104",
		X"11AB",
		X"122C",
		X"12D3",
		X"1354",
		X"13FB",
		X"147C",
		X"1523",
		X"15A4",
		X"164B",
		X"16CC",
		X"1773",
		X"17F4",
		X"189B",
		X"191C",
		X"19C3",
		X"1A44",
		X"1AEB",
		X"1B6C",
		X"1C13",
		X"1C94",
		X"1D3B",
		X"1DBC",
		X"1E63",
		X"1EE4",
		X"1F8B",
		X"200C",
		X"20B3",
		X"2134",
		X"21DB",
		X"225C",
		X"002B",
		X"00AC",
		X"0153",
		X"01D4",
		X"027B",
		X"02FC",
		X"03A3",
		X"0424",
		X"04CB",
		X"054C",
		X"05F3",
		X"0674",
		X"071B",
		X"079C",
		X"0843",
		X"08C4",
		X"096B",
		X"09EC",
		X"0A93",
		X"0B14",
		X"0BBB",
		X"0C3C",
		X"0CE3",
		X"0D64",
		X"0E0B",
		X"0E8C",
		X"0F33",
		X"0FB4",
		X"105B",
		X"10DC",
		X"1183",
		X"1204",
		X"12AB",
		X"132C",
		X"13D3",
		X"1454",
		X"14FB",
		X"157C",
		X"1623",
		X"16A4",
		X"174B",
		X"17CC",
		X"1873",
		X"18F4",
		X"199B",
		X"1A1C",
		X"1AC3",
		X"1B44",
		X"1BEB",
		X"1C6C",
		X"1D13",
		X"1D94",
		X"1E3B",
		X"1EBC",
		X"1F63",
		X"1FE4",
		X"208B",
		X"210C",
		X"21B3",
		X"2234",
		X"0003",
		X"0084",
		X"012B",
		X"01AC",
		X"0253",
		X"02D4",
		X"037B",
		X"03FC",
		X"04A3",
		X"0524",
		X"05CB",
		X"064C",
		X"06F3",
		X"0774",
		X"081B",
		X"089C",
		X"0943",
		X"09C4",
		X"0A6B",
		X"0AEC",
		X"0B93",
		X"0C14",
		X"0CBB",
		X"0D3C",
		X"0DE3",
		X"0E64",
		X"0F0B",
		X"0F8C",
		X"1033",
		X"10B4",
		X"115B",
		X"11DC",
		X"1283",
		X"1304",
		X"13AB",
		X"142C",
		X"14D3",
		X"1554",
		X"15FB",
		X"167C",
		X"1723",
		X"17A4",
		X"184B",
		X"18CC",
		X"1973",
		X"19F4",
		X"1A9B",
		X"1B1C",
		X"1BC3",
		X"1C44",
		X"1CEB",
		X"1D6C",
		X"1E13",
		X"1E94",
		X"1F3B",
		X"1FBC",
		X"2063",
		X"20E4",
		X"218B",
		X"220C",
		X"22B3",
		X"005C",
		X"0103",
		X"0184",
		X"022B",
		X"02AC",
		X"0353",
		X"03D4",
		X"047B",
		X"04FC",
		X"05A3",
		X"0624",
		X"06CB",
		X"074C",
		X"07F3",
		X"0874",
		X"091B",
		X"099C",
		X"0A43",
		X"0AC4",
		X"0B6B",
		X"0BEC",
		X"0C93",
		X"0D14",
		X"0DBB",
		X"0E3C",
		X"0EE3",
		X"0F64",
		X"100B",
		X"108C",
		X"1133",
		X"11B4",
		X"125B",
		X"12DC",
		X"1383",
		X"1404",
		X"14AB",
		X"152C",
		X"15D3",
		X"1654",
		X"16FB",
		X"177C",
		X"1823",
		X"18A4",
		X"194B",
		X"19CC",
		X"1A73",
		X"1AF4",
		X"1B9B",
		X"1C1C",
		X"1CC3",
		X"1D44",
		X"1DEB",
		X"1E6C",
		X"1F13",
		X"1F94",
		X"203B",
		X"20BC",
		X"2163",
		X"21E4",
		X"228B",
		X"0034",
		X"00DB",
		X"015C",
		X"0203",
		X"0284",
		X"032B",
		X"03AC",
		X"0453",
		X"04D4",
		X"057B",
		X"05FC",
		X"06A3",
		X"0724",
		X"07CB",
		X"084C",
		X"08F3",
		X"0974",
		X"0A1B",
		X"0A9C",
		X"0B43",
		X"0BC4",
		X"0C6B",
		X"0CEC",
		X"0D93",
		X"0E14",
		X"0EBB",
		X"0F3C",
		X"0FE3",
		X"1064",
		X"110B",
		X"118C",
		X"1233",
		X"12B4",
		X"135B",
		X"13DC",
		X"1483",
		X"1504",
		X"15AB",
		X"162C",
		X"16D3",
		X"1754",
		X"17FB",
		X"187C",
		X"1923",
		X"19A4",
		X"1A4B",
		X"1ACC",
		X"1B73",
		X"1BF4",
		X"1C9B",
		X"1D1C",
		X"1DC3",
		X"1E44",
		X"1EEB",
		X"1F6C",
		X"2013",
		X"2094",
		X"213B",
		X"21BC",
		X"2263",
		X"000C",
		X"00B3",
		X"0134",
		X"01DB",
		X"025C",
		X"0303",
		X"0384",
		X"042B",
		X"04AC",
		X"0553",
		X"05D4",
		X"067B",
		X"06FC",
		X"07A3",
		X"0824",
		X"08CB",
		X"094C",
		X"09F3",
		X"0A74",
		X"0B1B",
		X"0B9C",
		X"0C43",
		X"0CC4",
		X"0D6B",
		X"0DEC",
		X"0E93",
		X"0F14",
		X"0FBB",
		X"103C",
		X"10E3",
		X"1164",
		X"120B",
		X"128C",
		X"1333",
		X"13B4",
		X"145B",
		X"14DC",
		X"1583",
		X"1604",
		X"16AB",
		X"172C",
		X"17D3",
		X"1854",
		X"18FB",
		X"197C",
		X"1A23",
		X"1AA4",
		X"1B4B",
		X"1BCC",
		X"1C73",
		X"1CF4",
		X"1D9B",
		X"1E1C",
		X"1EC3",
		X"1F44",
		X"1FEB",
		X"206C",
		X"2113",
		X"2194",
		X"223B",
		X"22BC",
		X"008B",
		X"010C",
		X"01B3",
		X"0234",
		X"02DB",
		X"035C",
		X"0403",
		X"0484",
		X"052B",
		X"05AC",
		X"0653",
		X"06D4",
		X"077B",
		X"07FC",
		X"08A3",
		X"0924",
		X"09CB",
		X"0A4C",
		X"0AF3",
		X"0B74",
		X"0C1B",
		X"0C9C",
		X"0D43",
		X"0DC4",
		X"0E6B",
		X"0EEC",
		X"0F93",
		X"1014",
		X"10BB",
		X"113C",
		X"11E3",
		X"1264",
		X"130B",
		X"138C",
		X"1433",
		X"14B4",
		X"155B",
		X"15DC",
		X"1683",
		X"1704",
		X"17AB",
		X"182C",
		X"18D3",
		X"1954",
		X"19FB",
		X"1A7C",
		X"1B23",
		X"1BA4",
		X"1C4B",
		X"1CCC",
		X"1D73",
		X"1DF4",
		X"1E9B",
		X"1F1C",
		X"1FC3",
		X"2044",
		X"20EB",
		X"216C",
		X"2213",
		X"2294",
		X"0063",
		X"00E4",
		X"018B",
		X"020C",
		X"02B3",
		X"0334",
		X"03DB",
		X"045C",
		X"0503",
		X"0584",
		X"062B",
		X"06AC",
		X"0753",
		X"07D4",
		X"087B",
		X"08FC",
		X"09A3",
		X"0A24",
		X"0ACB",
		X"0B4C",
		X"0BF3",
		X"0C74",
		X"0D1B",
		X"0D9C",
		X"0E43",
		X"0EC4",
		X"0F6B",
		X"0FEC",
		X"1093",
		X"1114",
		X"11BB",
		X"123C",
		X"12E3",
		X"1364",
		X"140B",
		X"148C",
		X"1533",
		X"15B4",
		X"165B",
		X"16DC",
		X"1783",
		X"1804",
		X"18AB",
		X"192C",
		X"19D3",
		X"1A54",
		X"1AFB",
		X"1B7C",
		X"1C23",
		X"1CA4",
		X"1D4B",
		X"1DCC",
		X"1E73",
		X"1EF4",
		X"1F9B",
		X"201C",
		X"20C3",
		X"2144",
		X"21EB",
		X"226C",
		X"003B",
		X"00BC",
		X"0163",
		X"01E4",
		X"028B",
		X"030C",
		X"03B3",
		X"0434",
		X"04DB",
		X"055C",
		X"0603",
		X"0684",
		X"072B",
		X"07AC",
		X"0853",
		X"08D4",
		X"097B",
		X"09FC",
		X"0AA3",
		X"0B24",
		X"0BCB",
		X"0C4C",
		X"0CF3",
		X"0D74",
		X"0E1B",
		X"0E9C",
		X"0F43",
		X"0FC4",
		X"106B",
		X"10EC",
		X"1193",
		X"1214",
		X"12BB",
		X"133C",
		X"13E3",
		X"1464",
		X"150B",
		X"158C",
		X"1633",
		X"16B4",
		X"175B",
		X"17DC",
		X"1883",
		X"1904",
		X"19AB",
		X"1A2C",
		X"1AD3",
		X"1B54",
		X"1BFB",
		X"1C7C",
		X"1D23",
		X"1DA4",
		X"1E4B",
		X"1ECC",
		X"1F73",
		X"1FF4",
		X"209B",
		X"211C",
		X"21C3",
		X"2244",
		X"0013",
		X"0094",
		X"013B",
		X"01BC",
		X"0263",
		X"02E4",
		X"038B",
		X"040C",
		X"04B3",
		X"0534",
		X"05DB",
		X"065C",
		X"0703",
		X"0784",
		X"082B",
		X"08AC",
		X"0953",
		X"09D4",
		X"0A7B",
		X"0AFC",
		X"0BA3",
		X"0C24",
		X"0CCB",
		X"0D4C",
		X"0DF3",
		X"0E74",
		X"0F1B",
		X"0F9C",
		X"1043",
		X"10C4",
		X"116B",
		X"11EC",
		X"1293",
		X"1314",
		X"13BB",
		X"143C",
		X"14E3",
		X"1564",
		X"160B",
		X"168C",
		X"1733",
		X"17B4",
		X"185B",
		X"18DC",
		X"1983",
		X"1A04",
		X"1AAB",
		X"1B2C",
		X"1BD3",
		X"1C54",
		X"1CFB",
		X"1D7C",
		X"1E23",
		X"1EA4",
		X"1F4B",
		X"1FCC",
		X"2073",
		X"20F4",
		X"219B",
		X"221C",
		X"22C3",
		X"006C",
		X"0113",
		X"0194",
		X"023B",
		X"02BC",
		X"0363",
		X"03E4",
		X"048B",
		X"050C",
		X"05B3",
		X"0634",
		X"06DB",
		X"075C",
		X"0803",
		X"0884",
		X"092B",
		X"09AC",
		X"0A53",
		X"0AD4",
		X"0B7B",
		X"0BFC",
		X"0CA3",
		X"0D24",
		X"0DCB",
		X"0E4C",
		X"0EF3",
		X"0F74",
		X"101B",
		X"109C",
		X"1143",
		X"11C4",
		X"126B",
		X"12EC",
		X"1393",
		X"1414",
		X"14BB",
		X"153C",
		X"15E3",
		X"1664",
		X"170B",
		X"178C",
		X"1833",
		X"18B4",
		X"195B",
		X"19DC",
		X"1A83",
		X"1B04",
		X"1BAB",
		X"1C2C",
		X"1CD3",
		X"1D54",
		X"1DFB",
		X"1E7C",
		X"1F23",
		X"1FA4",
		X"204B",
		X"20CC",
		X"2173",
		X"21F4",
		X"229B",
		X"0044",
		X"00EB",
		X"016C",
		X"0213",
		X"0294",
		X"033B",
		X"03BC",
		X"0463",
		X"04E4",
		X"058B",
		X"060C",
		X"06B3",
		X"0734",
		X"07DB",
		X"085C",
		X"0903",
		X"0984",
		X"0A2B",
		X"0AAC",
		X"0B53",
		X"0BD4",
		X"0C7B",
		X"0CFC",
		X"0DA3",
		X"0E24",
		X"0ECB",
		X"0F4C",
		X"0FF3",
		X"1074",
		X"111B",
		X"119C",
		X"1243",
		X"12C4",
		X"136B",
		X"13EC",
		X"1493",
		X"1514",
		X"15BB",
		X"163C",
		X"16E3",
		X"1764",
		X"180B",
		X"188C",
		X"1933",
		X"19B4",
		X"1A5B",
		X"1ADC",
		X"1B83",
		X"1C04",
		X"1CAB",
		X"1D2C",
		X"1DD3",
		X"1E54",
		X"1EFB",
		X"1F7C",
		X"2023",
		X"20A4",
		X"214B",
		X"21CC",
		X"2273",
		X"001C",
		X"00C3",
		X"0144",
		X"01EB",
		X"026C",
		X"0313",
		X"0394",
		X"043B",
		X"04BC",
		X"0563",
		X"05E4",
		X"068B",
		X"070C",
		X"07B3",
		X"0834",
		X"08DB",
		X"095C",
		X"0A03",
		X"0A84",
		X"0B2B",
		X"0BAC",
		X"0C53",
		X"0CD4",
		X"0D7B",
		X"0DFC",
		X"0EA3",
		X"0F24",
		X"0FCB",
		X"104C",
		X"10F3",
		X"1174",
		X"121B",
		X"129C",
		X"1343",
		X"13C4",
		X"146B",
		X"14EC",
		X"1593",
		X"1614",
		X"16BB",
		X"173C",
		X"17E3",
		X"1864",
		X"190B",
		X"198C",
		X"1A33",
		X"1AB4",
		X"1B5B",
		X"1BDC",
		X"1C83",
		X"1D04",
		X"1DAB",
		X"1E2C",
		X"1ED3",
		X"1F54",
		X"1FFB",
		X"207C",
		X"2123",
		X"21A4",
		X"224B",
		X"22CC",
		X"009B",
		X"011C",
		X"01C3",
		X"0244",
		X"02EB",
		X"036C",
		X"0413",
		X"0494",
		X"053B",
		X"05BC",
		X"0663",
		X"06E4",
		X"078B",
		X"080C",
		X"08B3",
		X"0934",
		X"09DB",
		X"0A5C",
		X"0B03",
		X"0B84",
		X"0C2B",
		X"0CAC",
		X"0D53",
		X"0DD4",
		X"0E7B",
		X"0EFC",
		X"0FA3",
		X"1024",
		X"10CB",
		X"114C",
		X"11F3",
		X"1274",
		X"131B",
		X"139C",
		X"1443",
		X"14C4",
		X"156B",
		X"15EC",
		X"1693",
		X"1714",
		X"17BB",
		X"183C",
		X"18E3",
		X"1964",
		X"1A0B",
		X"1A8C",
		X"1B33",
		X"1BB4",
		X"1C5B",
		X"1CDC",
		X"1D83",
		X"1E04",
		X"1EAB",
		X"1F2C",
		X"1FD3",
		X"2054",
		X"20FB",
		X"217C",
		X"2223",
		X"22A4",
		X"0073",
		X"00F4",
		X"019B",
		X"021C",
		X"02C3",
		X"0344",
		X"03EB",
		X"046C",
		X"0513",
		X"0594",
		X"063B",
		X"06BC",
		X"0763",
		X"07E4",
		X"088B",
		X"090C",
		X"09B3",
		X"0A34",
		X"0ADB",
		X"0B5C",
		X"0C03",
		X"0C84",
		X"0D2B",
		X"0DAC",
		X"0E53",
		X"0ED4",
		X"0F7B",
		X"0FFC",
		X"10A3",
		X"1124",
		X"11CB",
		X"124C",
		X"12F3",
		X"1374",
		X"141B",
		X"149C",
		X"1543",
		X"15C4",
		X"166B",
		X"16EC",
		X"1793",
		X"1814",
		X"18BB",
		X"193C",
		X"19E3",
		X"1A64",
		X"1B0B",
		X"1B8C",
		X"1C33",
		X"1CB4",
		X"1D5B",
		X"1DDC",
		X"1E83",
		X"1F04",
		X"1FAB",
		X"202C",
		X"20D3",
		X"2154",
		X"21FB",
		X"227C",
		X"004B",
		X"00CC",
		X"0173",
		X"01F4",
		X"029B",
		X"031C",
		X"03C3",
		X"0444",
		X"04EB",
		X"056C",
		X"0613",
		X"0694",
		X"073B",
		X"07BC",
		X"0863",
		X"08E4",
		X"098B",
		X"0A0C",
		X"0AB3",
		X"0B34",
		X"0BDB",
		X"0C5C",
		X"0D03",
		X"0D84",
		X"0E2B",
		X"0EAC",
		X"0F53",
		X"0FD4",
		X"107B",
		X"10FC",
		X"11A3",
		X"1224",
		X"12CB",
		X"134C",
		X"13F3",
		X"1474",
		X"151B",
		X"159C",
		X"1643",
		X"16C4",
		X"176B",
		X"17EC",
		X"1893",
		X"1914",
		X"19BB",
		X"1A3C",
		X"1AE3",
		X"1B64",
		X"1C0B",
		X"1C8C",
		X"1D33",
		X"1DB4",
		X"1E5B",
		X"1EDC",
		X"1F83",
		X"2004",
		X"20AB",
		X"212C",
		X"21D3",
		X"2254",
		X"0023",
		X"00A4",
		X"014B",
		X"01CC",
		X"0273",
		X"02F4",
		X"039B",
		X"041C",
		X"04C3",
		X"0544",
		X"05EB",
		X"066C",
		X"0713",
		X"0794",
		X"083B",
		X"08BC",
		X"0963",
		X"09E4",
		X"0A8B",
		X"0B0C",
		X"0BB3",
		X"0C34",
		X"0CDB",
		X"0D5C",
		X"0E03",
		X"0E84",
		X"0F2B",
		X"0FAC",
		X"1053",
		X"10D4",
		X"117B",
		X"11FC",
		X"12A3",
		X"1324",
		X"13CB",
		X"144C",
		X"14F3",
		X"1574",
		X"161B",
		X"169C",
		X"1743",
		X"17C4",
		X"186B",
		X"18EC",
		X"1993",
		X"1A14",
		X"1ABB",
		X"1B3C",
		X"1BE3",
		X"1C64",
		X"1D0B",
		X"1D8C",
		X"1E33",
		X"1EB4",
		X"1F5B",
		X"1FDC",
		X"2083",
		X"2104",
		X"21AB",
		X"222C",
		X"22D3",
		X"007C",
		X"0123",
		X"01A4",
		X"024B",
		X"02CC",
		X"0373",
		X"03F4",
		X"049B",
		X"051C",
		X"05C3",
		X"0644",
		X"06EB",
		X"076C",
		X"0813",
		X"0894",
		X"093B",
		X"09BC",
		X"0A63",
		X"0AE4",
		X"0B8B",
		X"0C0C",
		X"0CB3",
		X"0D34",
		X"0DDB",
		X"0E5C",
		X"0F03",
		X"0F84",
		X"102B",
		X"10AC",
		X"1153",
		X"11D4",
		X"127B",
		X"12FC",
		X"13A3",
		X"1424",
		X"14CB",
		X"154C",
		X"15F3",
		X"1674",
		X"171B",
		X"179C",
		X"1843",
		X"18C4",
		X"196B",
		X"19EC",
		X"1A93",
		X"1B14",
		X"1BBB",
		X"1C3C",
		X"1CE3",
		X"1D64",
		X"1E0B",
		X"1E8C",
		X"1F33",
		X"1FB4",
		X"205B",
		X"20DC",
		X"2183",
		X"2204",
		X"22AB",
		X"0054",
		X"00FB",
		X"017C",
		X"0223",
		X"02A4",
		X"034B",
		X"03CC",
		X"0473",
		X"04F4",
		X"059B",
		X"061C",
		X"06C3",
		X"0744",
		X"07EB",
		X"086C",
		X"0913",
		X"0994",
		X"0A3B",
		X"0ABC",
		X"0B63",
		X"0BE4",
		X"0C8B",
		X"0D0C",
		X"0DB3",
		X"0E34",
		X"0EDB",
		X"0F5C",
		X"1003",
		X"1084",
		X"112B",
		X"11AC",
		X"1253",
		X"12D4",
		X"137B",
		X"13FC",
		X"14A3",
		X"1524",
		X"15CB",
		X"164C",
		X"16F3",
		X"1774",
		X"181B",
		X"189C",
		X"1943",
		X"19C4",
		X"1A6B",
		X"1AEC",
		X"1B93",
		X"1C14",
		X"1CBB",
		X"1D3C",
		X"1DE3",
		X"1E64",
		X"1F0B",
		X"1F8C",
		X"2033",
		X"20B4",
		X"215B",
		X"21DC",
		X"2283",
		X"002C",
		X"00D3",
		X"0154",
		X"01FB",
		X"027C",
		X"0323",
		X"03A4",
		X"044B",
		X"04CC",
		X"0573",
		X"05F4",
		X"069B",
		X"071C",
		X"07C3",
		X"0844",
		X"08EB",
		X"096C",
		X"0A13",
		X"0A94",
		X"0B3B",
		X"0BBC",
		X"0C63",
		X"0CE4",
		X"0D8B",
		X"0E0C",
		X"0EB3",
		X"0F34",
		X"0FDB",
		X"105C",
		X"1103",
		X"1184",
		X"122B",
		X"12AC",
		X"1353",
		X"13D4",
		X"147B",
		X"14FC",
		X"15A3",
		X"1624",
		X"16CB",
		X"174C",
		X"17F3",
		X"1874",
		X"191B",
		X"199C",
		X"1A43",
		X"1AC4",
		X"1B6B",
		X"1BEC",
		X"1C93",
		X"1D14",
		X"1DBB",
		X"1E3C",
		X"1EE3",
		X"1F64",
		X"200B",
		X"208C",
		X"2133",
		X"21B4",
		X"225B",
		X"0002",
		X"00A9",
		X"00FA",
		X"01A1",
		X"01F2",
		X"0299",
		X"02EA",
		X"0391",
		X"03E2",
		X"0489",
		X"04DA",
		X"0581",
		X"05D2",
		X"0679",
		X"06CA",
		X"0771",
		X"07C2",
		X"0869",
		X"08BA",
		X"0961",
		X"09B2",
		X"0A59",
		X"0AAA",
		X"0B51",
		X"0BA2",
		X"0C49",
		X"0C9A",
		X"0D41",
		X"0D92",
		X"0E39",
		X"0E8A",
		X"0F31",
		X"0F82",
		X"1029",
		X"107A",
		X"1121",
		X"1172",
		X"1219",
		X"126A",
		X"1311",
		X"1362",
		X"1409",
		X"145A",
		X"1501",
		X"1552",
		X"15F9",
		X"164A",
		X"16F1",
		X"1742",
		X"17E9",
		X"183A",
		X"18E1",
		X"1932",
		X"19D9",
		X"1A2A",
		X"1AD1",
		X"1B22",
		X"1BC9",
		X"1C1A",
		X"1CC1",
		X"1D12",
		X"1DB9",
		X"1E0A",
		X"1EB1",
		X"1F02",
		X"1FA9",
		X"1FFA",
		X"20A1",
		X"20F2",
		X"2199",
		X"21EA",
		X"2291",
		X"000A",
		X"00B1",
		X"0102",
		X"01A9",
		X"01FA",
		X"02A1",
		X"02F2",
		X"0399",
		X"03EA",
		X"0491",
		X"04E2",
		X"0589",
		X"05DA",
		X"0681",
		X"06D2",
		X"0779",
		X"07CA",
		X"0871",
		X"08C2",
		X"0969",
		X"09BA",
		X"0A61",
		X"0AB2",
		X"0B59",
		X"0BAA",
		X"0C51",
		X"0CA2",
		X"0D49",
		X"0D9A",
		X"0E41",
		X"0E92",
		X"0F39",
		X"0F8A",
		X"1031",
		X"1082",
		X"1129",
		X"117A",
		X"1221",
		X"1272",
		X"1319",
		X"136A",
		X"1411",
		X"1462",
		X"1509",
		X"155A",
		X"1601",
		X"1652",
		X"16F9",
		X"174A",
		X"17F1",
		X"1842",
		X"18E9",
		X"193A",
		X"19E1",
		X"1A32",
		X"1AD9",
		X"1B2A",
		X"1BD1",
		X"1C22",
		X"1CC9",
		X"1D1A",
		X"1DC1",
		X"1E12",
		X"1EB9",
		X"1F0A",
		X"1FB1",
		X"2002",
		X"20A9",
		X"20FA",
		X"21A1",
		X"21F2",
		X"2299",
		X"0012",
		X"00B9",
		X"010A",
		X"01B1",
		X"0202",
		X"02A9",
		X"02FA",
		X"03A1",
		X"03F2",
		X"0499",
		X"04EA",
		X"0591",
		X"05E2",
		X"0689",
		X"06DA",
		X"0781",
		X"07D2",
		X"0879",
		X"08CA",
		X"0971",
		X"09C2",
		X"0A69",
		X"0ABA",
		X"0B61",
		X"0BB2",
		X"0C59",
		X"0CAA",
		X"0D51",
		X"0DA2",
		X"0E49",
		X"0E9A",
		X"0F41",
		X"0F92",
		X"1039",
		X"108A",
		X"1131",
		X"1182",
		X"1229",
		X"127A",
		X"1321",
		X"1372",
		X"1419",
		X"146A",
		X"1511",
		X"1562",
		X"1609",
		X"165A",
		X"1701",
		X"1752",
		X"17F9",
		X"184A",
		X"18F1",
		X"1942",
		X"19E9",
		X"1A3A",
		X"1AE1",
		X"1B32",
		X"1BD9",
		X"1C2A",
		X"1CD1",
		X"1D22",
		X"1DC9",
		X"1E1A",
		X"1EC1",
		X"1F12",
		X"1FB9",
		X"200A",
		X"20B1",
		X"2102",
		X"21A9",
		X"21FA",
		X"22A1",
		X"001A",
		X"00C1",
		X"0112",
		X"01B9",
		X"020A",
		X"02B1",
		X"0302",
		X"03A9",
		X"03FA",
		X"04A1",
		X"04F2",
		X"0599",
		X"05EA",
		X"0691",
		X"06E2",
		X"0789",
		X"07DA",
		X"0881",
		X"08D2",
		X"0979",
		X"09CA",
		X"0A71",
		X"0AC2",
		X"0B69",
		X"0BBA",
		X"0C61",
		X"0CB2",
		X"0D59",
		X"0DAA",
		X"0E51",
		X"0EA2",
		X"0F49",
		X"0F9A",
		X"1041",
		X"1092",
		X"1139",
		X"118A",
		X"1231",
		X"1282",
		X"1329",
		X"137A",
		X"1421",
		X"1472",
		X"1519",
		X"156A",
		X"1611",
		X"1662",
		X"1709",
		X"175A",
		X"1801",
		X"1852",
		X"18F9",
		X"194A",
		X"19F1",
		X"1A42",
		X"1AE9",
		X"1B3A",
		X"1BE1",
		X"1C32",
		X"1CD9",
		X"1D2A",
		X"1DD1",
		X"1E22",
		X"1EC9",
		X"1F1A",
		X"1FC1",
		X"2012",
		X"20B9",
		X"210A",
		X"21B1",
		X"2202",
		X"22A9",
		X"0022",
		X"00C9",
		X"011A",
		X"01C1",
		X"0212",
		X"02B9",
		X"030A",
		X"03B1",
		X"0402",
		X"04A9",
		X"04FA",
		X"05A1",
		X"05F2",
		X"0699",
		X"06EA",
		X"0791",
		X"07E2",
		X"0889",
		X"08DA",
		X"0981",
		X"09D2",
		X"0A79",
		X"0ACA",
		X"0B71",
		X"0BC2",
		X"0C69",
		X"0CBA",
		X"0D61",
		X"0DB2",
		X"0E59",
		X"0EAA",
		X"0F51",
		X"0FA2",
		X"1049",
		X"109A",
		X"1141",
		X"1192",
		X"1239",
		X"128A",
		X"1331",
		X"1382",
		X"1429",
		X"147A",
		X"1521",
		X"1572",
		X"1619",
		X"166A",
		X"1711",
		X"1762",
		X"1809",
		X"185A",
		X"1901",
		X"1952",
		X"19F9",
		X"1A4A",
		X"1AF1",
		X"1B42",
		X"1BE9",
		X"1C3A",
		X"1CE1",
		X"1D32",
		X"1DD9",
		X"1E2A",
		X"1ED1",
		X"1F22",
		X"1FC9",
		X"201A",
		X"20C1",
		X"2112",
		X"21B9",
		X"220A",
		X"22B1",
		X"002A",
		X"00D1",
		X"0122",
		X"01C9",
		X"021A",
		X"02C1",
		X"0312",
		X"03B9",
		X"040A",
		X"04B1",
		X"0502",
		X"05A9",
		X"05FA",
		X"06A1",
		X"06F2",
		X"0799",
		X"07EA",
		X"0891",
		X"08E2",
		X"0989",
		X"09DA",
		X"0A81",
		X"0AD2",
		X"0B79",
		X"0BCA",
		X"0C71",
		X"0CC2",
		X"0D69",
		X"0DBA",
		X"0E61",
		X"0EB2",
		X"0F59",
		X"0FAA",
		X"1051",
		X"10A2",
		X"1149",
		X"119A",
		X"1241",
		X"1292",
		X"1339",
		X"138A",
		X"1431",
		X"1482",
		X"1529",
		X"157A",
		X"1621",
		X"1672",
		X"1719",
		X"176A",
		X"1811",
		X"1862",
		X"1909",
		X"195A",
		X"1A01",
		X"1A52",
		X"1AF9",
		X"1B4A",
		X"1BF1",
		X"1C42",
		X"1CE9",
		X"1D3A",
		X"1DE1",
		X"1E32",
		X"1ED9",
		X"1F2A",
		X"1FD1",
		X"2022",
		X"20C9",
		X"211A",
		X"21C1",
		X"2212",
		X"22B9",
		X"0032",
		X"00D9",
		X"012A",
		X"01D1",
		X"0222",
		X"02C9",
		X"031A",
		X"03C1",
		X"0412",
		X"04B9",
		X"050A",
		X"05B1",
		X"0602",
		X"06A9",
		X"06FA",
		X"07A1",
		X"07F2",
		X"0899",
		X"08EA",
		X"0991",
		X"09E2",
		X"0A89",
		X"0ADA",
		X"0B81",
		X"0BD2",
		X"0C79",
		X"0CCA",
		X"0D71",
		X"0DC2",
		X"0E69",
		X"0EBA",
		X"0F61",
		X"0FB2",
		X"1059",
		X"10AA",
		X"1151",
		X"11A2",
		X"1249",
		X"129A",
		X"1341",
		X"1392",
		X"1439",
		X"148A",
		X"1531",
		X"1582",
		X"1629",
		X"167A",
		X"1721",
		X"1772",
		X"1819",
		X"186A",
		X"1911",
		X"1962",
		X"1A09",
		X"1A5A",
		X"1B01",
		X"1B52",
		X"1BF9",
		X"1C4A",
		X"1CF1",
		X"1D42",
		X"1DE9",
		X"1E3A",
		X"1EE1",
		X"1F32",
		X"1FD9",
		X"202A",
		X"20D1",
		X"2122",
		X"21C9",
		X"221A",
		X"22C1",
		X"003A",
		X"00E1",
		X"0132",
		X"01D9",
		X"022A",
		X"02D1",
		X"0322",
		X"03C9",
		X"041A",
		X"04C1",
		X"0512",
		X"05B9",
		X"060A",
		X"06B1",
		X"0702",
		X"07A9",
		X"07FA",
		X"08A1",
		X"08F2",
		X"0999",
		X"09EA",
		X"0A91",
		X"0AE2",
		X"0B89",
		X"0BDA",
		X"0C81",
		X"0CD2",
		X"0D79",
		X"0DCA",
		X"0E71",
		X"0EC2",
		X"0F69",
		X"0FBA",
		X"1061",
		X"10B2",
		X"1159",
		X"11AA",
		X"1251",
		X"12A2",
		X"1349",
		X"139A",
		X"1441",
		X"1492",
		X"1539",
		X"158A",
		X"1631",
		X"1682",
		X"1729",
		X"177A",
		X"1821",
		X"1872",
		X"1919",
		X"196A",
		X"1A11",
		X"1A62",
		X"1B09",
		X"1B5A",
		X"1C01",
		X"1C52",
		X"1CF9",
		X"1D4A",
		X"1DF1",
		X"1E42",
		X"1EE9",
		X"1F3A",
		X"1FE1",
		X"2032",
		X"20D9",
		X"212A",
		X"21D1",
		X"2222",
		X"22C9",
		X"0042",
		X"00E9",
		X"013A",
		X"01E1",
		X"0232",
		X"02D9",
		X"032A",
		X"03D1",
		X"0422",
		X"04C9",
		X"051A",
		X"05C1",
		X"0612",
		X"06B9",
		X"070A",
		X"07B1",
		X"0802",
		X"08A9",
		X"08FA",
		X"09A1",
		X"09F2",
		X"0A99",
		X"0AEA",
		X"0B91",
		X"0BE2",
		X"0C89",
		X"0CDA",
		X"0D81",
		X"0DD2",
		X"0E79",
		X"0ECA",
		X"0F71",
		X"0FC2",
		X"1069",
		X"10BA",
		X"1161",
		X"11B2",
		X"1259",
		X"12AA",
		X"1351",
		X"13A2",
		X"1449",
		X"149A",
		X"1541",
		X"1592",
		X"1639",
		X"168A",
		X"1731",
		X"1782",
		X"1829",
		X"187A",
		X"1921",
		X"1972",
		X"1A19",
		X"1A6A",
		X"1B11",
		X"1B62",
		X"1C09",
		X"1C5A",
		X"1D01",
		X"1D52",
		X"1DF9",
		X"1E4A",
		X"1EF1",
		X"1F42",
		X"1FE9",
		X"203A",
		X"20E1",
		X"2132",
		X"21D9",
		X"222A",
		X"22D1",
		X"004A",
		X"00F1",
		X"0142",
		X"01E9",
		X"023A",
		X"02E1",
		X"0332",
		X"03D9",
		X"042A",
		X"04D1",
		X"0522",
		X"05C9",
		X"061A",
		X"06C1",
		X"0712",
		X"07B9",
		X"080A",
		X"08B1",
		X"0902",
		X"09A9",
		X"09FA",
		X"0AA1",
		X"0AF2",
		X"0B99",
		X"0BEA",
		X"0C91",
		X"0CE2",
		X"0D89",
		X"0DDA",
		X"0E81",
		X"0ED2",
		X"0F79",
		X"0FCA",
		X"1071",
		X"10C2",
		X"1169",
		X"11BA",
		X"1261",
		X"12B2",
		X"1359",
		X"13AA",
		X"1451",
		X"14A2",
		X"1549",
		X"159A",
		X"1641",
		X"1692",
		X"1739",
		X"178A",
		X"1831",
		X"1882",
		X"1929",
		X"197A",
		X"1A21",
		X"1A72",
		X"1B19",
		X"1B6A",
		X"1C11",
		X"1C62",
		X"1D09",
		X"1D5A",
		X"1E01",
		X"1E52",
		X"1EF9",
		X"1F4A",
		X"1FF1",
		X"2042",
		X"20E9",
		X"213A",
		X"21E1",
		X"2232",
		X"0001",
		X"0052",
		X"00F9",
		X"014A",
		X"01F1",
		X"0242",
		X"02E9",
		X"033A",
		X"03E1",
		X"0432",
		X"04D9",
		X"052A",
		X"05D1",
		X"0622",
		X"06C9",
		X"071A",
		X"07C1",
		X"0812",
		X"08B9",
		X"090A",
		X"09B1",
		X"0A02",
		X"0AA9",
		X"0AFA",
		X"0BA1",
		X"0BF2",
		X"0C99",
		X"0CEA",
		X"0D91",
		X"0DE2",
		X"0E89",
		X"0EDA",
		X"0F81",
		X"0FD2",
		X"1079",
		X"10CA",
		X"1171",
		X"11C2",
		X"1269",
		X"12BA",
		X"1361",
		X"13B2",
		X"1459",
		X"14AA",
		X"1551",
		X"15A2",
		X"1649",
		X"169A",
		X"1741",
		X"1792",
		X"1839",
		X"188A",
		X"1931",
		X"1982",
		X"1A29",
		X"1A7A",
		X"1B21",
		X"1B72",
		X"1C19",
		X"1C6A",
		X"1D11",
		X"1D62",
		X"1E09",
		X"1E5A",
		X"1F01",
		X"1F52",
		X"1FF9",
		X"204A",
		X"20F1",
		X"2142",
		X"21E9",
		X"223A",
		X"0009",
		X"005A",
		X"0101",
		X"0152",
		X"01F9",
		X"024A",
		X"02F1",
		X"0342",
		X"03E9",
		X"043A",
		X"04E1",
		X"0532",
		X"05D9",
		X"062A",
		X"06D1",
		X"0722",
		X"07C9",
		X"081A",
		X"08C1",
		X"0912",
		X"09B9",
		X"0A0A",
		X"0AB1",
		X"0B02",
		X"0BA9",
		X"0BFA",
		X"0CA1",
		X"0CF2",
		X"0D99",
		X"0DEA",
		X"0E91",
		X"0EE2",
		X"0F89",
		X"0FDA",
		X"1081",
		X"10D2",
		X"1179",
		X"11CA",
		X"1271",
		X"12C2",
		X"1369",
		X"13BA",
		X"1461",
		X"14B2",
		X"1559",
		X"15AA",
		X"1651",
		X"16A2",
		X"1749",
		X"179A",
		X"1841",
		X"1892",
		X"1939",
		X"198A",
		X"1A31",
		X"1A82",
		X"1B29",
		X"1B7A",
		X"1C21",
		X"1C72",
		X"1D19",
		X"1D6A",
		X"1E11",
		X"1E62",
		X"1F09",
		X"1F5A",
		X"2001",
		X"2052",
		X"20F9",
		X"214A",
		X"21F1",
		X"2242",
		X"0011",
		X"0062",
		X"0109",
		X"015A",
		X"0201",
		X"0252",
		X"02F9",
		X"034A",
		X"03F1",
		X"0442",
		X"04E9",
		X"053A",
		X"05E1",
		X"0632",
		X"06D9",
		X"072A",
		X"07D1",
		X"0822",
		X"08C9",
		X"091A",
		X"09C1",
		X"0A12",
		X"0AB9",
		X"0B0A",
		X"0BB1",
		X"0C02",
		X"0CA9",
		X"0CFA",
		X"0DA1",
		X"0DF2",
		X"0E99",
		X"0EEA",
		X"0F91",
		X"0FE2",
		X"1089",
		X"10DA",
		X"1181",
		X"11D2",
		X"1279",
		X"12CA",
		X"1371",
		X"13C2",
		X"1469",
		X"14BA",
		X"1561",
		X"15B2",
		X"1659",
		X"16AA",
		X"1751",
		X"17A2",
		X"1849",
		X"189A",
		X"1941",
		X"1992",
		X"1A39",
		X"1A8A",
		X"1B31",
		X"1B82",
		X"1C29",
		X"1C7A",
		X"1D21",
		X"1D72",
		X"1E19",
		X"1E6A",
		X"1F11",
		X"1F62",
		X"2009",
		X"205A",
		X"2101",
		X"2152",
		X"21F9",
		X"224A",
		X"0019",
		X"006A",
		X"0111",
		X"0162",
		X"0209",
		X"025A",
		X"0301",
		X"0352",
		X"03F9",
		X"044A",
		X"04F1",
		X"0542",
		X"05E9",
		X"063A",
		X"06E1",
		X"0732",
		X"07D9",
		X"082A",
		X"08D1",
		X"0922",
		X"09C9",
		X"0A1A",
		X"0AC1",
		X"0B12",
		X"0BB9",
		X"0C0A",
		X"0CB1",
		X"0D02",
		X"0DA9",
		X"0DFA",
		X"0EA1",
		X"0EF2",
		X"0F99",
		X"0FEA",
		X"1091",
		X"10E2",
		X"1189",
		X"11DA",
		X"1281",
		X"12D2",
		X"1379",
		X"13CA",
		X"1471",
		X"14C2",
		X"1569",
		X"15BA",
		X"1661",
		X"16B2",
		X"1759",
		X"17AA",
		X"1851",
		X"18A2",
		X"1949",
		X"199A",
		X"1A41",
		X"1A92",
		X"1B39",
		X"1B8A",
		X"1C31",
		X"1C82",
		X"1D29",
		X"1D7A",
		X"1E21",
		X"1E72",
		X"1F19",
		X"1F6A",
		X"2011",
		X"2062",
		X"2109",
		X"215A",
		X"2201",
		X"2252",
		X"0021",
		X"0072",
		X"0119",
		X"016A",
		X"0211",
		X"0262",
		X"0309",
		X"035A",
		X"0401",
		X"0452",
		X"04F9",
		X"054A",
		X"05F1",
		X"0642",
		X"06E9",
		X"073A",
		X"07E1",
		X"0832",
		X"08D9",
		X"092A",
		X"09D1",
		X"0A22",
		X"0AC9",
		X"0B1A",
		X"0BC1",
		X"0C12",
		X"0CB9",
		X"0D0A",
		X"0DB1",
		X"0E02",
		X"0EA9",
		X"0EFA",
		X"0FA1",
		X"0FF2",
		X"1099",
		X"10EA",
		X"1191",
		X"11E2",
		X"1289",
		X"12DA",
		X"1381",
		X"13D2",
		X"1479",
		X"14CA",
		X"1571",
		X"15C2",
		X"1669",
		X"16BA",
		X"1761",
		X"17B2",
		X"1859",
		X"18AA",
		X"1951",
		X"19A2",
		X"1A49",
		X"1A9A",
		X"1B41",
		X"1B92",
		X"1C39",
		X"1C8A",
		X"1D31",
		X"1D82",
		X"1E29",
		X"1E7A",
		X"1F21",
		X"1F72",
		X"2019",
		X"206A",
		X"2111",
		X"2162",
		X"2209",
		X"225A",
		X"0029",
		X"007A",
		X"0121",
		X"0172",
		X"0219",
		X"026A",
		X"0311",
		X"0362",
		X"0409",
		X"045A",
		X"0501",
		X"0552",
		X"05F9",
		X"064A",
		X"06F1",
		X"0742",
		X"07E9",
		X"083A",
		X"08E1",
		X"0932",
		X"09D9",
		X"0A2A",
		X"0AD1",
		X"0B22",
		X"0BC9",
		X"0C1A",
		X"0CC1",
		X"0D12",
		X"0DB9",
		X"0E0A",
		X"0EB1",
		X"0F02",
		X"0FA9",
		X"0FFA",
		X"10A1",
		X"10F2",
		X"1199",
		X"11EA",
		X"1291",
		X"12E2",
		X"1389",
		X"13DA",
		X"1481",
		X"14D2",
		X"1579",
		X"15CA",
		X"1671",
		X"16C2",
		X"1769",
		X"17BA",
		X"1861",
		X"18B2",
		X"1959",
		X"19AA",
		X"1A51",
		X"1AA2",
		X"1B49",
		X"1B9A",
		X"1C41",
		X"1C92",
		X"1D39",
		X"1D8A",
		X"1E31",
		X"1E82",
		X"1F29",
		X"1F7A",
		X"2021",
		X"2072",
		X"2119",
		X"216A",
		X"2211",
		X"2262",
		X"0031",
		X"0082",
		X"0129",
		X"017A",
		X"0221",
		X"0272",
		X"0319",
		X"036A",
		X"0411",
		X"0462",
		X"0509",
		X"055A",
		X"0601",
		X"0652",
		X"06F9",
		X"074A",
		X"07F1",
		X"0842",
		X"08E9",
		X"093A",
		X"09E1",
		X"0A32",
		X"0AD9",
		X"0B2A",
		X"0BD1",
		X"0C22",
		X"0CC9",
		X"0D1A",
		X"0DC1",
		X"0E12",
		X"0EB9",
		X"0F0A",
		X"0FB1",
		X"1002",
		X"10A9",
		X"10FA",
		X"11A1",
		X"11F2",
		X"1299",
		X"12EA",
		X"1391",
		X"13E2",
		X"1489",
		X"14DA",
		X"1581",
		X"15D2",
		X"1679",
		X"16CA",
		X"1771",
		X"17C2",
		X"1869",
		X"18BA",
		X"1961",
		X"19B2",
		X"1A59",
		X"1AAA",
		X"1B51",
		X"1BA2",
		X"1C49",
		X"1C9A",
		X"1D41",
		X"1D92",
		X"1E39",
		X"1E8A",
		X"1F31",
		X"1F82",
		X"2029",
		X"207A",
		X"2121",
		X"2172",
		X"2219",
		X"226A",
		X"0039",
		X"008A",
		X"0131",
		X"0182",
		X"0229",
		X"027A",
		X"0321",
		X"0372",
		X"0419",
		X"046A",
		X"0511",
		X"0562",
		X"0609",
		X"065A",
		X"0701",
		X"0752",
		X"07F9",
		X"084A",
		X"08F1",
		X"0942",
		X"09E9",
		X"0A3A",
		X"0AE1",
		X"0B32",
		X"0BD9",
		X"0C2A",
		X"0CD1",
		X"0D22",
		X"0DC9",
		X"0E1A",
		X"0EC1",
		X"0F12",
		X"0FB9",
		X"100A",
		X"10B1",
		X"1102",
		X"11A9",
		X"11FA",
		X"12A1",
		X"12F2",
		X"1399",
		X"13EA",
		X"1491",
		X"14E2",
		X"1589",
		X"15DA",
		X"1681",
		X"16D2",
		X"1779",
		X"17CA",
		X"1871",
		X"18C2",
		X"1969",
		X"19BA",
		X"1A61",
		X"1AB2",
		X"1B59",
		X"1BAA",
		X"1C51",
		X"1CA2",
		X"1D49",
		X"1D9A",
		X"1E41",
		X"1E92",
		X"1F39",
		X"1F8A",
		X"2031",
		X"2082",
		X"2129",
		X"217A",
		X"2221",
		X"2272",
		X"0041",
		X"0092",
		X"0139",
		X"018A",
		X"0231",
		X"0282",
		X"0329",
		X"037A",
		X"0421",
		X"0472",
		X"0519",
		X"056A",
		X"0611",
		X"0662",
		X"0709",
		X"075A",
		X"0801",
		X"0852",
		X"08F9",
		X"094A",
		X"09F1",
		X"0A42",
		X"0AE9",
		X"0B3A",
		X"0BE1",
		X"0C32",
		X"0CD9",
		X"0D2A",
		X"0DD1",
		X"0E22",
		X"0EC9",
		X"0F1A",
		X"0FC1",
		X"1012",
		X"10B9",
		X"110A",
		X"11B1",
		X"1202",
		X"12A9",
		X"12FA",
		X"13A1",
		X"13F2",
		X"1499",
		X"14EA",
		X"1591",
		X"15E2",
		X"1689",
		X"16DA",
		X"1781",
		X"17D2",
		X"1879",
		X"18CA",
		X"1971",
		X"19C2",
		X"1A69",
		X"1ABA",
		X"1B61",
		X"1BB2",
		X"1C59",
		X"1CAA",
		X"1D51",
		X"1DA2",
		X"1E49",
		X"1E9A",
		X"1F41",
		X"1F92",
		X"2039",
		X"208A",
		X"2131",
		X"2182",
		X"2229",
		X"227A",
		X"0049",
		X"009A",
		X"0141",
		X"0192",
		X"0239",
		X"028A",
		X"0331",
		X"0382",
		X"0429",
		X"047A",
		X"0521",
		X"0572",
		X"0619",
		X"066A",
		X"0711",
		X"0762",
		X"0809",
		X"085A",
		X"0901",
		X"0952",
		X"09F9",
		X"0A4A",
		X"0AF1",
		X"0B42",
		X"0BE9",
		X"0C3A",
		X"0CE1",
		X"0D32",
		X"0DD9",
		X"0E2A",
		X"0ED1",
		X"0F22",
		X"0FC9",
		X"101A",
		X"10C1",
		X"1112",
		X"11B9",
		X"120A",
		X"12B1",
		X"1302",
		X"13A9",
		X"13FA",
		X"14A1",
		X"14F2",
		X"1599",
		X"15EA",
		X"1691",
		X"16E2",
		X"1789",
		X"17DA",
		X"1881",
		X"18D2",
		X"1979",
		X"19CA",
		X"1A71",
		X"1AC2",
		X"1B69",
		X"1BBA",
		X"1C61",
		X"1CB2",
		X"1D59",
		X"1DAA",
		X"1E51",
		X"1EA2",
		X"1F49",
		X"1F9A",
		X"2041",
		X"2092",
		X"2139",
		X"218A",
		X"2231",
		X"2282",
		X"0051",
		X"00A2",
		X"0149",
		X"019A",
		X"0241",
		X"0292",
		X"0339",
		X"038A",
		X"0431",
		X"0482",
		X"0529",
		X"057A",
		X"0621",
		X"0672",
		X"0719",
		X"076A",
		X"0811",
		X"0862",
		X"0909",
		X"095A",
		X"0A01",
		X"0A52",
		X"0AF9",
		X"0B4A",
		X"0BF1",
		X"0C42",
		X"0CE9",
		X"0D3A",
		X"0DE1",
		X"0E32",
		X"0ED9",
		X"0F2A",
		X"0FD1",
		X"1022",
		X"10C9",
		X"111A",
		X"11C1",
		X"1212",
		X"12B9",
		X"130A",
		X"13B1",
		X"1402",
		X"14A9",
		X"14FA",
		X"15A1",
		X"15F2",
		X"1699",
		X"16EA",
		X"1791",
		X"17E2",
		X"1889",
		X"18DA",
		X"1981",
		X"19D2",
		X"1A79",
		X"1ACA",
		X"1B71",
		X"1BC2",
		X"1C69",
		X"1CBA",
		X"1D61",
		X"1DB2",
		X"1E59",
		X"1EAA",
		X"1F51",
		X"1FA2",
		X"2049",
		X"209A",
		X"2141",
		X"2192",
		X"2239",
		X"228A",
		X"0059",
		X"00AA",
		X"0151",
		X"01A2",
		X"0249",
		X"029A",
		X"0341",
		X"0392",
		X"0439",
		X"048A",
		X"0531",
		X"0582",
		X"0629",
		X"067A",
		X"0721",
		X"0772",
		X"0819",
		X"086A",
		X"0911",
		X"0962",
		X"0A09",
		X"0A5A",
		X"0B01",
		X"0B52",
		X"0BF9",
		X"0C4A",
		X"0CF1",
		X"0D42",
		X"0DE9",
		X"0E3A",
		X"0EE1",
		X"0F32",
		X"0FD9",
		X"102A",
		X"10D1",
		X"1122",
		X"11C9",
		X"121A",
		X"12C1",
		X"1312",
		X"13B9",
		X"140A",
		X"14B1",
		X"1502",
		X"15A9",
		X"15FA",
		X"16A1",
		X"16F2",
		X"1799",
		X"17EA",
		X"1891",
		X"18E2",
		X"1989",
		X"19DA",
		X"1A81",
		X"1AD2",
		X"1B79",
		X"1BCA",
		X"1C71",
		X"1CC2",
		X"1D69",
		X"1DBA",
		X"1E61",
		X"1EB2",
		X"1F59",
		X"1FAA",
		X"2051",
		X"20A2",
		X"2149",
		X"219A",
		X"2241",
		X"2292",
		X"0061",
		X"00B2",
		X"0159",
		X"01AA",
		X"0251",
		X"02A2",
		X"0349",
		X"039A",
		X"0441",
		X"0492",
		X"0539",
		X"058A",
		X"0631",
		X"0682",
		X"0729",
		X"077A",
		X"0821",
		X"0872",
		X"0919",
		X"096A",
		X"0A11",
		X"0A62",
		X"0B09",
		X"0B5A",
		X"0C01",
		X"0C52",
		X"0CF9",
		X"0D4A",
		X"0DF1",
		X"0E42",
		X"0EE9",
		X"0F3A",
		X"0FE1",
		X"1032",
		X"10D9",
		X"112A",
		X"11D1",
		X"1222",
		X"12C9",
		X"131A",
		X"13C1",
		X"1412",
		X"14B9",
		X"150A",
		X"15B1",
		X"1602",
		X"16A9",
		X"16FA",
		X"17A1",
		X"17F2",
		X"1899",
		X"18EA",
		X"1991",
		X"19E2",
		X"1A89",
		X"1ADA",
		X"1B81",
		X"1BD2",
		X"1C79",
		X"1CCA",
		X"1D71",
		X"1DC2",
		X"1E69",
		X"1EBA",
		X"1F61",
		X"1FB2",
		X"2059",
		X"20AA",
		X"2151",
		X"21A2",
		X"2249",
		X"229A",
		X"0069",
		X"00BA",
		X"0161",
		X"01B2",
		X"0259",
		X"02AA",
		X"0351",
		X"03A2",
		X"0449",
		X"049A",
		X"0541",
		X"0592",
		X"0639",
		X"068A",
		X"0731",
		X"0782",
		X"0829",
		X"087A",
		X"0921",
		X"0972",
		X"0A19",
		X"0A6A",
		X"0B11",
		X"0B62",
		X"0C09",
		X"0C5A",
		X"0D01",
		X"0D52",
		X"0DF9",
		X"0E4A",
		X"0EF1",
		X"0F42",
		X"0FE9",
		X"103A",
		X"10E1",
		X"1132",
		X"11D9",
		X"122A",
		X"12D1",
		X"1322",
		X"13C9",
		X"141A",
		X"14C1",
		X"1512",
		X"15B9",
		X"160A",
		X"16B1",
		X"1702",
		X"17A9",
		X"17FA",
		X"18A1",
		X"18F2",
		X"1999",
		X"19EA",
		X"1A91",
		X"1AE2",
		X"1B89",
		X"1BDA",
		X"1C81",
		X"1CD2",
		X"1D79",
		X"1DCA",
		X"1E71",
		X"1EC2",
		X"1F69",
		X"1FBA",
		X"2061",
		X"20B2",
		X"2159",
		X"21AA",
		X"2251",
		X"22A2",
		X"0071",
		X"00C2",
		X"0169",
		X"01BA",
		X"0261",
		X"02B2",
		X"0359",
		X"03AA",
		X"0451",
		X"04A2",
		X"0549",
		X"059A",
		X"0641",
		X"0692",
		X"0739",
		X"078A",
		X"0831",
		X"0882",
		X"0929",
		X"097A",
		X"0A21",
		X"0A72",
		X"0B19",
		X"0B6A",
		X"0C11",
		X"0C62",
		X"0D09",
		X"0D5A",
		X"0E01",
		X"0E52",
		X"0EF9",
		X"0F4A",
		X"0FF1",
		X"1042",
		X"10E9",
		X"113A",
		X"11E1",
		X"1232",
		X"12D9",
		X"132A",
		X"13D1",
		X"1422",
		X"14C9",
		X"151A",
		X"15C1",
		X"1612",
		X"16B9",
		X"170A",
		X"17B1",
		X"1802",
		X"18A9",
		X"18FA",
		X"19A1",
		X"19F2",
		X"1A99",
		X"1AEA",
		X"1B91",
		X"1BE2",
		X"1C89",
		X"1CDA",
		X"1D81",
		X"1DD2",
		X"1E79",
		X"1ECA",
		X"1F71",
		X"1FC2",
		X"2069",
		X"20BA",
		X"2161",
		X"21B2",
		X"2259",
		X"22AA",
		X"0079",
		X"00CA",
		X"0171",
		X"01C2",
		X"0269",
		X"02BA",
		X"0361",
		X"03B2",
		X"0459",
		X"04AA",
		X"0551",
		X"05A2",
		X"0649",
		X"069A",
		X"0741",
		X"0792",
		X"0839",
		X"088A",
		X"0931",
		X"0982",
		X"0A29",
		X"0A7A",
		X"0B21",
		X"0B72",
		X"0C19",
		X"0C6A",
		X"0D11",
		X"0D62",
		X"0E09",
		X"0E5A",
		X"0F01",
		X"0F52",
		X"0FF9",
		X"104A",
		X"10F1",
		X"1142",
		X"11E9",
		X"123A",
		X"12E1",
		X"1332",
		X"13D9",
		X"142A",
		X"14D1",
		X"1522",
		X"15C9",
		X"161A",
		X"16C1",
		X"1712",
		X"17B9",
		X"180A",
		X"18B1",
		X"1902",
		X"19A9",
		X"19FA",
		X"1AA1",
		X"1AF2",
		X"1B99",
		X"1BEA",
		X"1C91",
		X"1CE2",
		X"1D89",
		X"1DDA",
		X"1E81",
		X"1ED2",
		X"1F79",
		X"1FCA",
		X"2071",
		X"20C2",
		X"2169",
		X"21BA",
		X"2261",
		X"22B2",
		X"0081",
		X"00D2",
		X"0179",
		X"01CA",
		X"0271",
		X"02C2",
		X"0369",
		X"03BA",
		X"0461",
		X"04B2",
		X"0559",
		X"05AA",
		X"0651",
		X"06A2",
		X"0749",
		X"079A",
		X"0841",
		X"0892",
		X"0939",
		X"098A",
		X"0A31",
		X"0A82",
		X"0B29",
		X"0B7A",
		X"0C21",
		X"0C72",
		X"0D19",
		X"0D6A",
		X"0E11",
		X"0E62",
		X"0F09",
		X"0F5A",
		X"1001",
		X"1052",
		X"10F9",
		X"114A",
		X"11F1",
		X"1242",
		X"12E9",
		X"133A",
		X"13E1",
		X"1432",
		X"14D9",
		X"152A",
		X"15D1",
		X"1622",
		X"16C9",
		X"171A",
		X"17C1",
		X"1812",
		X"18B9",
		X"190A",
		X"19B1",
		X"1A02",
		X"1AA9",
		X"1AFA",
		X"1BA1",
		X"1BF2",
		X"1C99",
		X"1CEA",
		X"1D91",
		X"1DE2",
		X"1E89",
		X"1EDA",
		X"1F81",
		X"1FD2",
		X"2079",
		X"20CA",
		X"2171",
		X"21C2",
		X"2269",
		X"22BA",
		X"0089",
		X"00DA",
		X"0181",
		X"01D2",
		X"0279",
		X"02CA",
		X"0371",
		X"03C2",
		X"0469",
		X"04BA",
		X"0561",
		X"05B2",
		X"0659",
		X"06AA",
		X"0751",
		X"07A2",
		X"0849",
		X"089A",
		X"0941",
		X"0992",
		X"0A39",
		X"0A8A",
		X"0B31",
		X"0B82",
		X"0C29",
		X"0C7A",
		X"0D21",
		X"0D72",
		X"0E19",
		X"0E6A",
		X"0F11",
		X"0F62",
		X"1009",
		X"105A",
		X"1101",
		X"1152",
		X"11F9",
		X"124A",
		X"12F1",
		X"1342",
		X"13E9",
		X"143A",
		X"14E1",
		X"1532",
		X"15D9",
		X"162A",
		X"16D1",
		X"1722",
		X"17C9",
		X"181A",
		X"18C1",
		X"1912",
		X"19B9",
		X"1A0A",
		X"1AB1",
		X"1B02",
		X"1BA9",
		X"1BFA",
		X"1CA1",
		X"1CF2",
		X"1D99",
		X"1DEA",
		X"1E91",
		X"1EE2",
		X"1F89",
		X"1FDA",
		X"2081",
		X"20D2",
		X"2179",
		X"21CA",
		X"2271",
		X"22C2",
		X"0091",
		X"00E2",
		X"0189",
		X"01DA",
		X"0281",
		X"02D2",
		X"0379",
		X"03CA",
		X"0471",
		X"04C2",
		X"0569",
		X"05BA",
		X"0661",
		X"06B2",
		X"0759",
		X"07AA",
		X"0851",
		X"08A2",
		X"0949",
		X"099A",
		X"0A41",
		X"0A92",
		X"0B39",
		X"0B8A",
		X"0C31",
		X"0C82",
		X"0D29",
		X"0D7A",
		X"0E21",
		X"0E72",
		X"0F19",
		X"0F6A",
		X"1011",
		X"1062",
		X"1109",
		X"115A",
		X"1201",
		X"1252",
		X"12F9",
		X"134A",
		X"13F1",
		X"1442",
		X"14E9",
		X"153A",
		X"15E1",
		X"1632",
		X"16D9",
		X"172A",
		X"17D1",
		X"1822",
		X"18C9",
		X"191A",
		X"19C1",
		X"1A12",
		X"1AB9",
		X"1B0A",
		X"1BB1",
		X"1C02",
		X"1CA9",
		X"1CFA",
		X"1DA1",
		X"1DF2",
		X"1E99",
		X"1EEA",
		X"1F91",
		X"1FE2",
		X"2089",
		X"20DA",
		X"2181",
		X"21D2",
		X"2279",
		X"22CA",
		X"0099",
		X"00EA",
		X"0191",
		X"01E2",
		X"0289",
		X"02DA",
		X"0381",
		X"03D2",
		X"0479",
		X"04CA",
		X"0571",
		X"05C2",
		X"0669",
		X"06BA",
		X"0761",
		X"07B2",
		X"0859",
		X"08AA",
		X"0951",
		X"09A2",
		X"0A49",
		X"0A9A",
		X"0B41",
		X"0B92",
		X"0C39",
		X"0C8A",
		X"0D31",
		X"0D82",
		X"0E29",
		X"0E7A",
		X"0F21",
		X"0F72",
		X"1019",
		X"106A",
		X"1111",
		X"1162",
		X"1209",
		X"125A",
		X"1301",
		X"1352",
		X"13F9",
		X"144A",
		X"14F1",
		X"1542",
		X"15E9",
		X"163A",
		X"16E1",
		X"1732",
		X"17D9",
		X"182A",
		X"18D1",
		X"1922",
		X"19C9",
		X"1A1A",
		X"1AC1",
		X"1B12",
		X"1BB9",
		X"1C0A",
		X"1CB1",
		X"1D02",
		X"1DA9",
		X"1DFA",
		X"1EA1",
		X"1EF2",
		X"1F99",
		X"1FEA",
		X"2091",
		X"20E2",
		X"2189",
		X"21DA",
		X"2281",
		X"22D2",
		X"00A1",
		X"00F2",
		X"0199",
		X"01EA",
		X"0291",
		X"02E2",
		X"0389",
		X"03DA",
		X"0481",
		X"04D2",
		X"0579",
		X"05CA",
		X"0671",
		X"06C2",
		X"0769",
		X"07BA",
		X"0861",
		X"08B2",
		X"0959",
		X"09AA",
		X"0A51",
		X"0AA2",
		X"0B49",
		X"0B9A",
		X"0C41",
		X"0C92",
		X"0D39",
		X"0D8A",
		X"0E31",
		X"0E82",
		X"0F29",
		X"0F7A",
		X"1021",
		X"1072",
		X"1119",
		X"116A",
		X"1211",
		X"1262",
		X"1309",
		X"135A",
		X"1401",
		X"1452",
		X"14F9",
		X"154A",
		X"15F1",
		X"1642",
		X"16E9",
		X"173A",
		X"17E1",
		X"1832",
		X"18D9",
		X"192A",
		X"19D1",
		X"1A22",
		X"1AC9",
		X"1B1A",
		X"1BC1",
		X"1C12",
		X"1CB9",
		X"1D0A",
		X"1DB1",
		X"1E02",
		X"1EA9",
		X"1EFA",
		X"1FA1",
		X"1FF2",
		X"2099",
		X"20EA",
		X"2191",
		X"21E2",
		X"2289",
		X"0008",
		X"00AF",
		X"0180",
		X"0227",
		X"02F8",
		X"039F",
		X"0470",
		X"0517",
		X"05E8",
		X"068F",
		X"0760",
		X"0807",
		X"08D8",
		X"097F",
		X"0A50",
		X"0AF7",
		X"0BC8",
		X"0C6F",
		X"0D40",
		X"0DE7",
		X"0EB8",
		X"0F5F",
		X"1030",
		X"10D7",
		X"11A8",
		X"124F",
		X"1320",
		X"13C7",
		X"1498",
		X"153F",
		X"1610",
		X"16B7",
		X"1788",
		X"182F",
		X"1900",
		X"19A7",
		X"1A78",
		X"1B1F",
		X"1BF0",
		X"1C97",
		X"1D68",
		X"1E0F",
		X"1EE0",
		X"1F87",
		X"2058",
		X"20FF",
		X"21D0",
		X"2277",
		X"0070",
		X"0117",
		X"01E8",
		X"028F",
		X"0360",
		X"0407",
		X"04D8",
		X"057F",
		X"0650",
		X"06F7",
		X"07C8",
		X"086F",
		X"0940",
		X"09E7",
		X"0AB8",
		X"0B5F",
		X"0C30",
		X"0CD7",
		X"0DA8",
		X"0E4F",
		X"0F20",
		X"0FC7",
		X"1098",
		X"113F",
		X"1210",
		X"12B7",
		X"1388",
		X"142F",
		X"1500",
		X"15A7",
		X"1678",
		X"171F",
		X"17F0",
		X"1897",
		X"1968",
		X"1A0F",
		X"1AE0",
		X"1B87",
		X"1C58",
		X"1CFF",
		X"1DD0",
		X"1E77",
		X"1F48",
		X"1FEF",
		X"20C0",
		X"2167",
		X"2238",
		X"0007",
		X"00D8",
		X"017F",
		X"0250",
		X"02F7",
		X"03C8",
		X"046F",
		X"0540",
		X"05E7",
		X"06B8",
		X"075F",
		X"0830",
		X"08D7",
		X"09A8",
		X"0A4F",
		X"0B20",
		X"0BC7",
		X"0C98",
		X"0D3F",
		X"0E10",
		X"0EB7",
		X"0F88",
		X"102F",
		X"1100",
		X"11A7",
		X"1278",
		X"131F",
		X"13F0",
		X"1497",
		X"1568",
		X"160F",
		X"16E0",
		X"1787",
		X"1858",
		X"18FF",
		X"19D0",
		X"1A77",
		X"1B48",
		X"1BEF",
		X"1CC0",
		X"1D67",
		X"1E38",
		X"1EDF",
		X"1FB0",
		X"2057",
		X"2128",
		X"21CF",
		X"22A0",
		X"006F",
		X"0140",
		X"01E7",
		X"02B8",
		X"035F",
		X"0430",
		X"04D7",
		X"05A8",
		X"064F",
		X"0720",
		X"07C7",
		X"0898",
		X"093F",
		X"0A10",
		X"0AB7",
		X"0B88",
		X"0C2F",
		X"0D00",
		X"0DA7",
		X"0E78",
		X"0F1F",
		X"0FF0",
		X"1097",
		X"1168",
		X"120F",
		X"12E0",
		X"1387",
		X"1458",
		X"14FF",
		X"15D0",
		X"1677",
		X"1748",
		X"17EF",
		X"18C0",
		X"1967",
		X"1A38",
		X"1ADF",
		X"1BB0",
		X"1C57",
		X"1D28",
		X"1DCF",
		X"1EA0",
		X"1F47",
		X"2018",
		X"20BF",
		X"2190",
		X"2237",
		X"0030",
		X"00D7",
		X"01A8",
		X"024F",
		X"0320",
		X"03C7",
		X"0498",
		X"053F",
		X"0610",
		X"06B7",
		X"0788",
		X"082F",
		X"0900",
		X"09A7",
		X"0A78",
		X"0B1F",
		X"0BF0",
		X"0C97",
		X"0D68",
		X"0E0F",
		X"0EE0",
		X"0F87",
		X"1058",
		X"10FF",
		X"11D0",
		X"1277",
		X"1348",
		X"13EF",
		X"14C0",
		X"1567",
		X"1638",
		X"16DF",
		X"17B0",
		X"1857",
		X"1928",
		X"19CF",
		X"1AA0",
		X"1B47",
		X"1C18",
		X"1CBF",
		X"1D90",
		X"1E37",
		X"1F08",
		X"1FAF",
		X"2080",
		X"2127",
		X"21F8",
		X"229F",
		X"0098",
		X"013F",
		X"0210",
		X"02B7",
		X"0388",
		X"042F",
		X"0500",
		X"05A7",
		X"0678",
		X"071F",
		X"07F0",
		X"0897",
		X"0968",
		X"0A0F",
		X"0AE0",
		X"0B87",
		X"0C58",
		X"0CFF",
		X"0DD0",
		X"0E77",
		X"0F48",
		X"0FEF",
		X"10C0",
		X"1167",
		X"1238",
		X"12DF",
		X"13B0",
		X"1457",
		X"1528",
		X"15CF",
		X"16A0",
		X"1747",
		X"1818",
		X"18BF",
		X"1990",
		X"1A37",
		X"1B08",
		X"1BAF",
		X"1C80",
		X"1D27",
		X"1DF8",
		X"1E9F",
		X"1F70",
		X"2017",
		X"20E8",
		X"218F",
		X"2260",
		X"002F",
		X"0100",
		X"01A7",
		X"0278",
		X"031F",
		X"03F0",
		X"0497",
		X"0568",
		X"060F",
		X"06E0",
		X"0787",
		X"0858",
		X"08FF",
		X"09D0",
		X"0A77",
		X"0B48",
		X"0BEF",
		X"0CC0",
		X"0D67",
		X"0E38",
		X"0EDF",
		X"0FB0",
		X"1057",
		X"1128",
		X"11CF",
		X"12A0",
		X"1347",
		X"1418",
		X"14BF",
		X"1590",
		X"1637",
		X"1708",
		X"17AF",
		X"1880",
		X"1927",
		X"19F8",
		X"1A9F",
		X"1B70",
		X"1C17",
		X"1CE8",
		X"1D8F",
		X"1E60",
		X"1F07",
		X"1FD8",
		X"207F",
		X"2150",
		X"21F7",
		X"22C8",
		X"0097",
		X"0168",
		X"020F",
		X"02E0",
		X"0387",
		X"0458",
		X"04FF",
		X"05D0",
		X"0677",
		X"0748",
		X"07EF",
		X"08C0",
		X"0967",
		X"0A38",
		X"0ADF",
		X"0BB0",
		X"0C57",
		X"0D28",
		X"0DCF",
		X"0EA0",
		X"0F47",
		X"1018",
		X"10BF",
		X"1190",
		X"1237",
		X"1308",
		X"13AF",
		X"1480",
		X"1527",
		X"15F8",
		X"169F",
		X"1770",
		X"1817",
		X"18E8",
		X"198F",
		X"1A60",
		X"1B07",
		X"1BD8",
		X"1C7F",
		X"1D50",
		X"1DF7",
		X"1EC8",
		X"1F6F",
		X"2040",
		X"20E7",
		X"21B8",
		X"225F",
		X"0058",
		X"00FF",
		X"01D0",
		X"0277",
		X"0348",
		X"03EF",
		X"04C0",
		X"0567",
		X"0638",
		X"06DF",
		X"07B0",
		X"0857",
		X"0928",
		X"09CF",
		X"0AA0",
		X"0B47",
		X"0C18",
		X"0CBF",
		X"0D90",
		X"0E37",
		X"0F08",
		X"0FAF",
		X"1080",
		X"1127",
		X"11F8",
		X"129F",
		X"1370",
		X"1417",
		X"14E8",
		X"158F",
		X"1660",
		X"1707",
		X"17D8",
		X"187F",
		X"1950",
		X"19F7",
		X"1AC8",
		X"1B6F",
		X"1C40",
		X"1CE7",
		X"1DB8",
		X"1E5F",
		X"1F30",
		X"1FD7",
		X"20A8",
		X"214F",
		X"2220",
		X"22C7",
		X"00C0",
		X"0167",
		X"0238",
		X"02DF",
		X"03B0",
		X"0457",
		X"0528",
		X"05CF",
		X"06A0",
		X"0747",
		X"0818",
		X"08BF",
		X"0990",
		X"0A37",
		X"0B08",
		X"0BAF",
		X"0C80",
		X"0D27",
		X"0DF8",
		X"0E9F",
		X"0F70",
		X"1017",
		X"10E8",
		X"118F",
		X"1260",
		X"1307",
		X"13D8",
		X"147F",
		X"1550",
		X"15F7",
		X"16C8",
		X"176F",
		X"1840",
		X"18E7",
		X"19B8",
		X"1A5F",
		X"1B30",
		X"1BD7",
		X"1CA8",
		X"1D4F",
		X"1E20",
		X"1EC7",
		X"1F98",
		X"203F",
		X"2110",
		X"21B7",
		X"2288",
		X"0057",
		X"0128",
		X"01CF",
		X"02A0",
		X"0347",
		X"0418",
		X"04BF",
		X"0590",
		X"0637",
		X"0708",
		X"07AF",
		X"0880",
		X"0927",
		X"09F8",
		X"0A9F",
		X"0B70",
		X"0C17",
		X"0CE8",
		X"0D8F",
		X"0E60",
		X"0F07",
		X"0FD8",
		X"107F",
		X"1150",
		X"11F7",
		X"12C8",
		X"136F",
		X"1440",
		X"14E7",
		X"15B8",
		X"165F",
		X"1730",
		X"17D7",
		X"18A8",
		X"194F",
		X"1A20",
		X"1AC7",
		X"1B98",
		X"1C3F",
		X"1D10",
		X"1DB7",
		X"1E88",
		X"1F2F",
		X"2000",
		X"20A7",
		X"2178",
		X"221F",
		X"0018",
		X"00BF",
		X"0190",
		X"0237",
		X"0308",
		X"03AF",
		X"0480",
		X"0527",
		X"05F8",
		X"069F",
		X"0770",
		X"0817",
		X"08E8",
		X"098F",
		X"0A60",
		X"0B07",
		X"0BD8",
		X"0C7F",
		X"0D50",
		X"0DF7",
		X"0EC8",
		X"0F6F",
		X"1040",
		X"10E7",
		X"11B8",
		X"125F",
		X"1330",
		X"13D7",
		X"14A8",
		X"154F",
		X"1620",
		X"16C7",
		X"1798",
		X"183F",
		X"1910",
		X"19B7",
		X"1A88",
		X"1B2F",
		X"1C00",
		X"1CA7",
		X"1D78",
		X"1E1F",
		X"1EF0",
		X"1F97",
		X"2068",
		X"210F",
		X"21E0",
		X"2287",
		X"0080",
		X"0127",
		X"01F8",
		X"029F",
		X"0370",
		X"0417",
		X"04E8",
		X"058F",
		X"0660",
		X"0707",
		X"07D8",
		X"087F",
		X"0950",
		X"09F7",
		X"0AC8",
		X"0B6F",
		X"0C40",
		X"0CE7",
		X"0DB8",
		X"0E5F",
		X"0F30",
		X"0FD7",
		X"10A8",
		X"114F",
		X"1220",
		X"12C7",
		X"1398",
		X"143F",
		X"1510",
		X"15B7",
		X"1688",
		X"172F",
		X"1800",
		X"18A7",
		X"1978",
		X"1A1F",
		X"1AF0",
		X"1B97",
		X"1C68",
		X"1D0F",
		X"1DE0",
		X"1E87",
		X"1F58",
		X"1FFF",
		X"20D0",
		X"2177",
		X"2248",
		X"0017",
		X"00E8",
		X"018F",
		X"0260",
		X"0307",
		X"03D8",
		X"047F",
		X"0550",
		X"05F7",
		X"06C8",
		X"076F",
		X"0840",
		X"08E7",
		X"09B8",
		X"0A5F",
		X"0B30",
		X"0BD7",
		X"0CA8",
		X"0D4F",
		X"0E20",
		X"0EC7",
		X"0F98",
		X"103F",
		X"1110",
		X"11B7",
		X"1288",
		X"132F",
		X"1400",
		X"14A7",
		X"1578",
		X"161F",
		X"16F0",
		X"1797",
		X"1868",
		X"190F",
		X"19E0",
		X"1A87",
		X"1B58",
		X"1BFF",
		X"1CD0",
		X"1D77",
		X"1E48",
		X"1EEF",
		X"1FC0",
		X"2067",
		X"2138",
		X"21DF",
		X"22B0",
		X"007F",
		X"0150",
		X"01F7",
		X"02C8",
		X"036F",
		X"0440",
		X"04E7",
		X"05B8",
		X"065F",
		X"0730",
		X"07D7",
		X"08A8",
		X"094F",
		X"0A20",
		X"0AC7",
		X"0B98",
		X"0C3F",
		X"0D10",
		X"0DB7",
		X"0E88",
		X"0F2F",
		X"1000",
		X"10A7",
		X"1178",
		X"121F",
		X"12F0",
		X"1397",
		X"1468",
		X"150F",
		X"15E0",
		X"1687",
		X"1758",
		X"17FF",
		X"18D0",
		X"1977",
		X"1A48",
		X"1AEF",
		X"1BC0",
		X"1C67",
		X"1D38",
		X"1DDF",
		X"1EB0",
		X"1F57",
		X"2028",
		X"20CF",
		X"21A0",
		X"2247",
		X"0040",
		X"00E7",
		X"01B8",
		X"025F",
		X"0330",
		X"03D7",
		X"04A8",
		X"054F",
		X"0620",
		X"06C7",
		X"0798",
		X"083F",
		X"0910",
		X"09B7",
		X"0A88",
		X"0B2F",
		X"0C00",
		X"0CA7",
		X"0D78",
		X"0E1F",
		X"0EF0",
		X"0F97",
		X"1068",
		X"110F",
		X"11E0",
		X"1287",
		X"1358",
		X"13FF",
		X"14D0",
		X"1577",
		X"1648",
		X"16EF",
		X"17C0",
		X"1867",
		X"1938",
		X"19DF",
		X"1AB0",
		X"1B57",
		X"1C28",
		X"1CCF",
		X"1DA0",
		X"1E47",
		X"1F18",
		X"1FBF",
		X"2090",
		X"2137",
		X"2208",
		X"22AF",
		X"00A8",
		X"014F",
		X"0220",
		X"02C7",
		X"0398",
		X"043F",
		X"0510",
		X"05B7",
		X"0688",
		X"072F",
		X"0800",
		X"08A7",
		X"0978",
		X"0A1F",
		X"0AF0",
		X"0B97",
		X"0C68",
		X"0D0F",
		X"0DE0",
		X"0E87",
		X"0F58",
		X"0FFF",
		X"10D0",
		X"1177",
		X"1248",
		X"12EF",
		X"13C0",
		X"1467",
		X"1538",
		X"15DF",
		X"16B0",
		X"1757",
		X"1828",
		X"18CF",
		X"19A0",
		X"1A47",
		X"1B18",
		X"1BBF",
		X"1C90",
		X"1D37",
		X"1E08",
		X"1EAF",
		X"1F80",
		X"2027",
		X"20F8",
		X"219F",
		X"2270",
		X"003F",
		X"0110",
		X"01B7",
		X"0288",
		X"032F",
		X"0400",
		X"04A7",
		X"0578",
		X"061F",
		X"06F0",
		X"0797",
		X"0868",
		X"090F",
		X"09E0",
		X"0A87",
		X"0B58",
		X"0BFF",
		X"0CD0",
		X"0D77",
		X"0E48",
		X"0EEF",
		X"0FC0",
		X"1067",
		X"1138",
		X"11DF",
		X"12B0",
		X"1357",
		X"1428",
		X"14CF",
		X"15A0",
		X"1647",
		X"1718",
		X"17BF",
		X"1890",
		X"1937",
		X"1A08",
		X"1AAF",
		X"1B80",
		X"1C27",
		X"1CF8",
		X"1D9F",
		X"1E70",
		X"1F17",
		X"1FE8",
		X"208F",
		X"2160",
		X"2207",
		X"22D8",
		X"00A7",
		X"0178",
		X"021F",
		X"02F0",
		X"0397",
		X"0468",
		X"050F",
		X"05E0",
		X"0687",
		X"0758",
		X"07FF",
		X"08D0",
		X"0977",
		X"0A48",
		X"0AEF",
		X"0BC0",
		X"0C67",
		X"0D38",
		X"0DDF",
		X"0EB0",
		X"0F57",
		X"1028",
		X"10CF",
		X"11A0",
		X"1247",
		X"1318",
		X"13BF",
		X"1490",
		X"1537",
		X"1608",
		X"16AF",
		X"1780",
		X"1827",
		X"18F8",
		X"199F",
		X"1A70",
		X"1B17",
		X"1BE8",
		X"1C8F",
		X"1D60",
		X"1E07",
		X"1ED8",
		X"1F7F",
		X"2050",
		X"20F7",
		X"21C8",
		X"226F",
		X"0068",
		X"010F",
		X"01E0",
		X"0287",
		X"0358",
		X"03FF",
		X"04D0",
		X"0577",
		X"0648",
		X"06EF",
		X"07C0",
		X"0867",
		X"0938",
		X"09DF",
		X"0AB0",
		X"0B57",
		X"0C28",
		X"0CCF",
		X"0DA0",
		X"0E47",
		X"0F18",
		X"0FBF",
		X"1090",
		X"1137",
		X"1208",
		X"12AF",
		X"1380",
		X"1427",
		X"14F8",
		X"159F",
		X"1670",
		X"1717",
		X"17E8",
		X"188F",
		X"1960",
		X"1A07",
		X"1AD8",
		X"1B7F",
		X"1C50",
		X"1CF7",
		X"1DC8",
		X"1E6F",
		X"1F40",
		X"1FE7",
		X"20B8",
		X"215F",
		X"2230",
		X"22D7",
		X"00D0",
		X"0177",
		X"0248",
		X"02EF",
		X"03C0",
		X"0467",
		X"0538",
		X"05DF",
		X"06B0",
		X"0757",
		X"0828",
		X"08CF",
		X"09A0",
		X"0A47",
		X"0B18",
		X"0BBF",
		X"0C90",
		X"0D37",
		X"0E08",
		X"0EAF",
		X"0F80",
		X"1027",
		X"10F8",
		X"119F",
		X"1270",
		X"1317",
		X"13E8",
		X"148F",
		X"1560",
		X"1607",
		X"16D8",
		X"177F",
		X"1850",
		X"18F7",
		X"19C8",
		X"1A6F",
		X"1B40",
		X"1BE7",
		X"1CB8",
		X"1D5F",
		X"1E30",
		X"1ED7",
		X"1FA8",
		X"204F",
		X"2120",
		X"21C7",
		X"2298",
		X"0067",
		X"0138",
		X"01DF",
		X"02B0",
		X"0357",
		X"0428",
		X"04CF",
		X"05A0",
		X"0647",
		X"0718",
		X"07BF",
		X"0890",
		X"0937",
		X"0A08",
		X"0AAF",
		X"0B80",
		X"0C27",
		X"0CF8",
		X"0D9F",
		X"0E70",
		X"0F17",
		X"0FE8",
		X"108F",
		X"1160",
		X"1207",
		X"12D8",
		X"137F",
		X"1450",
		X"14F7",
		X"15C8",
		X"166F",
		X"1740",
		X"17E7",
		X"18B8",
		X"195F",
		X"1A30",
		X"1AD7",
		X"1BA8",
		X"1C4F",
		X"1D20",
		X"1DC7",
		X"1E98",
		X"1F3F",
		X"2010",
		X"20B7",
		X"2188",
		X"222F",
		X"0028",
		X"00CF",
		X"01A0",
		X"0247",
		X"0318",
		X"03BF",
		X"0490",
		X"0537",
		X"0608",
		X"06AF",
		X"0780",
		X"0827",
		X"08F8",
		X"099F",
		X"0A70",
		X"0B17",
		X"0BE8",
		X"0C8F",
		X"0D60",
		X"0E07",
		X"0ED8",
		X"0F7F",
		X"1050",
		X"10F7",
		X"11C8",
		X"126F",
		X"1340",
		X"13E7",
		X"14B8",
		X"155F",
		X"1630",
		X"16D7",
		X"17A8",
		X"184F",
		X"1920",
		X"19C7",
		X"1A98",
		X"1B3F",
		X"1C10",
		X"1CB7",
		X"1D88",
		X"1E2F",
		X"1F00",
		X"1FA7",
		X"2078",
		X"211F",
		X"21F0",
		X"2297",
		X"0090",
		X"0137",
		X"0208",
		X"02AF",
		X"0380",
		X"0427",
		X"04F8",
		X"059F",
		X"0670",
		X"0717",
		X"07E8",
		X"088F",
		X"0960",
		X"0A07",
		X"0AD8",
		X"0B7F",
		X"0C50",
		X"0CF7",
		X"0DC8",
		X"0E6F",
		X"0F40",
		X"0FE7",
		X"10B8",
		X"115F",
		X"1230",
		X"12D7",
		X"13A8",
		X"144F",
		X"1520",
		X"15C7",
		X"1698",
		X"173F",
		X"1810",
		X"18B7",
		X"1988",
		X"1A2F",
		X"1B00",
		X"1BA7",
		X"1C78",
		X"1D1F",
		X"1DF0",
		X"1E97",
		X"1F68",
		X"200F",
		X"20E0",
		X"2187",
		X"2258",
		X"0027",
		X"00F8",
		X"019F",
		X"0270",
		X"0317",
		X"03E8",
		X"048F",
		X"0560",
		X"0607",
		X"06D8",
		X"077F",
		X"0850",
		X"08F7",
		X"09C8",
		X"0A6F",
		X"0B40",
		X"0BE7",
		X"0CB8",
		X"0D5F",
		X"0E30",
		X"0ED7",
		X"0FA8",
		X"104F",
		X"1120",
		X"11C7",
		X"1298",
		X"133F",
		X"1410",
		X"14B7",
		X"1588",
		X"162F",
		X"1700",
		X"17A7",
		X"1878",
		X"191F",
		X"19F0",
		X"1A97",
		X"1B68",
		X"1C0F",
		X"1CE0",
		X"1D87",
		X"1E58",
		X"1EFF",
		X"1FD0",
		X"2077",
		X"2148",
		X"21EF",
		X"22C0",
		X"008F",
		X"0160",
		X"0207",
		X"02D8",
		X"037F",
		X"0450",
		X"04F7",
		X"05C8",
		X"066F",
		X"0740",
		X"07E7",
		X"08B8",
		X"095F",
		X"0A30",
		X"0AD7",
		X"0BA8",
		X"0C4F",
		X"0D20",
		X"0DC7",
		X"0E98",
		X"0F3F",
		X"1010",
		X"10B7",
		X"1188",
		X"122F",
		X"1300",
		X"13A7",
		X"1478",
		X"151F",
		X"15F0",
		X"1697",
		X"1768",
		X"180F",
		X"18E0",
		X"1987",
		X"1A58",
		X"1AFF",
		X"1BD0",
		X"1C77",
		X"1D48",
		X"1DEF",
		X"1EC0",
		X"1F67",
		X"2038",
		X"20DF",
		X"21B0",
		X"2257",
		X"0050",
		X"00F7",
		X"01C8",
		X"026F",
		X"0340",
		X"03E7",
		X"04B8",
		X"055F",
		X"0630",
		X"06D7",
		X"07A8",
		X"084F",
		X"0920",
		X"09C7",
		X"0A98",
		X"0B3F",
		X"0C10",
		X"0CB7",
		X"0D88",
		X"0E2F",
		X"0F00",
		X"0FA7",
		X"1078",
		X"111F",
		X"11F0",
		X"1297",
		X"1368",
		X"140F",
		X"14E0",
		X"1587",
		X"1658",
		X"16FF",
		X"17D0",
		X"1877",
		X"1948",
		X"19EF",
		X"1AC0",
		X"1B67",
		X"1C38",
		X"1CDF",
		X"1DB0",
		X"1E57",
		X"1F28",
		X"1FCF",
		X"20A0",
		X"2147",
		X"2218",
		X"22BF",
		X"00B8",
		X"015F",
		X"0230",
		X"02D7",
		X"03A8",
		X"044F",
		X"0520",
		X"05C7",
		X"0698",
		X"073F",
		X"0810",
		X"08B7",
		X"0988",
		X"0A2F",
		X"0B00",
		X"0BA7",
		X"0C78",
		X"0D1F",
		X"0DF0",
		X"0E97",
		X"0F68",
		X"100F",
		X"10E0",
		X"1187",
		X"1258",
		X"12FF",
		X"13D0",
		X"1477",
		X"1548",
		X"15EF",
		X"16C0",
		X"1767",
		X"1838",
		X"18DF",
		X"19B0",
		X"1A57",
		X"1B28",
		X"1BCF",
		X"1CA0",
		X"1D47",
		X"1E18",
		X"1EBF",
		X"1F90",
		X"2037",
		X"2108",
		X"21AF",
		X"2280",
		X"004F",
		X"0120",
		X"01C7",
		X"0298",
		X"033F",
		X"0410",
		X"04B7",
		X"0588",
		X"062F",
		X"0700",
		X"07A7",
		X"0878",
		X"091F",
		X"09F0",
		X"0A97",
		X"0B68",
		X"0C0F",
		X"0CE0",
		X"0D87",
		X"0E58",
		X"0EFF",
		X"0FD0",
		X"1077",
		X"1148",
		X"11EF",
		X"12C0",
		X"1367",
		X"1438",
		X"14DF",
		X"15B0",
		X"1657",
		X"1728",
		X"17CF",
		X"18A0",
		X"1947",
		X"1A18",
		X"1ABF",
		X"1B90",
		X"1C37",
		X"1D08",
		X"1DAF",
		X"1E80",
		X"1F27",
		X"1FF8",
		X"209F",
		X"2170",
		X"2217",
		X"0010",
		X"00B7",
		X"0188",
		X"022F",
		X"0300",
		X"03A7",
		X"0478",
		X"051F",
		X"05F0",
		X"0697",
		X"0768",
		X"080F",
		X"08E0",
		X"0987",
		X"0A58",
		X"0AFF",
		X"0BD0",
		X"0C77",
		X"0D48",
		X"0DEF",
		X"0EC0",
		X"0F67",
		X"1038",
		X"10DF",
		X"11B0",
		X"1257",
		X"1328",
		X"13CF",
		X"14A0",
		X"1547",
		X"1618",
		X"16BF",
		X"1790",
		X"1837",
		X"1908",
		X"19AF",
		X"1A80",
		X"1B27",
		X"1BF8",
		X"1C9F",
		X"1D70",
		X"1E17",
		X"1EE8",
		X"1F8F",
		X"2060",
		X"2107",
		X"21D8",
		X"227F",
		X"0078",
		X"011F",
		X"01F0",
		X"0297",
		X"0368",
		X"040F",
		X"04E0",
		X"0587",
		X"0658",
		X"06FF",
		X"07D0",
		X"0877",
		X"0948",
		X"09EF",
		X"0AC0",
		X"0B67",
		X"0C38",
		X"0CDF",
		X"0DB0",
		X"0E57",
		X"0F28",
		X"0FCF",
		X"10A0",
		X"1147",
		X"1218",
		X"12BF",
		X"1390",
		X"1437",
		X"1508",
		X"15AF",
		X"1680",
		X"1727",
		X"17F8",
		X"189F",
		X"1970",
		X"1A17",
		X"1AE8",
		X"1B8F",
		X"1C60",
		X"1D07",
		X"1DD8",
		X"1E7F",
		X"1F50",
		X"1FF7",
		X"20C8",
		X"216F",
		X"2240",
		X"000F",
		X"00E0",
		X"0187",
		X"0258",
		X"02FF",
		X"03D0",
		X"0477",
		X"0548",
		X"05EF",
		X"06C0",
		X"0767",
		X"0838",
		X"08DF",
		X"09B0",
		X"0A57",
		X"0B28",
		X"0BCF",
		X"0CA0",
		X"0D47",
		X"0E18",
		X"0EBF",
		X"0F90",
		X"1037",
		X"1108",
		X"11AF",
		X"1280",
		X"1327",
		X"13F8",
		X"149F",
		X"1570",
		X"1617",
		X"16E8",
		X"178F",
		X"1860",
		X"1907",
		X"19D8",
		X"1A7F",
		X"1B50",
		X"1BF7",
		X"1CC8",
		X"1D6F",
		X"1E40",
		X"1EE7",
		X"1FB8",
		X"205F",
		X"2130",
		X"21D7",
		X"22A8",
		X"0077",
		X"0148",
		X"01EF",
		X"02C0",
		X"0367",
		X"0438",
		X"04DF",
		X"05B0",
		X"0657",
		X"0728",
		X"07CF",
		X"08A0",
		X"0947",
		X"0A18",
		X"0ABF",
		X"0B90",
		X"0C37",
		X"0D08",
		X"0DAF",
		X"0E80",
		X"0F27",
		X"0FF8",
		X"109F",
		X"1170",
		X"1217",
		X"12E8",
		X"138F",
		X"1460",
		X"1507",
		X"15D8",
		X"167F",
		X"1750",
		X"17F7",
		X"18C8",
		X"196F",
		X"1A40",
		X"1AE7",
		X"1BB8",
		X"1C5F",
		X"1D30",
		X"1DD7",
		X"1EA8",
		X"1F4F",
		X"2020",
		X"20C7",
		X"2198",
		X"223F",
		X"0038",
		X"00DF",
		X"01B0",
		X"0257",
		X"0328",
		X"03CF",
		X"04A0",
		X"0547",
		X"0618",
		X"06BF",
		X"0790",
		X"0837",
		X"0908",
		X"09AF",
		X"0A80",
		X"0B27",
		X"0BF8",
		X"0C9F",
		X"0D70",
		X"0E17",
		X"0EE8",
		X"0F8F",
		X"1060",
		X"1107",
		X"11D8",
		X"127F",
		X"1350",
		X"13F7",
		X"14C8",
		X"156F",
		X"1640",
		X"16E7",
		X"17B8",
		X"185F",
		X"1930",
		X"19D7",
		X"1AA8",
		X"1B4F",
		X"1C20",
		X"1CC7",
		X"1D98",
		X"1E3F",
		X"1F10",
		X"1FB7",
		X"2088",
		X"212F",
		X"2200",
		X"22A7",
		X"00A0",
		X"0147",
		X"0218",
		X"02BF",
		X"0390",
		X"0437",
		X"0508",
		X"05AF",
		X"0680",
		X"0727",
		X"07F8",
		X"089F",
		X"0970",
		X"0A17",
		X"0AE8",
		X"0B8F",
		X"0C60",
		X"0D07",
		X"0DD8",
		X"0E7F",
		X"0F50",
		X"0FF7",
		X"10C8",
		X"116F",
		X"1240",
		X"12E7",
		X"13B8",
		X"145F",
		X"1530",
		X"15D7",
		X"16A8",
		X"174F",
		X"1820",
		X"18C7",
		X"1998",
		X"1A3F",
		X"1B10",
		X"1BB7",
		X"1C88",
		X"1D2F",
		X"1E00",
		X"1EA7",
		X"1F78",
		X"201F",
		X"20F0",
		X"2197",
		X"2268",
		X"0037",
		X"0108",
		X"01AF",
		X"0280",
		X"0327",
		X"03F8",
		X"049F",
		X"0570",
		X"0617",
		X"06E8",
		X"078F",
		X"0860",
		X"0907",
		X"09D8",
		X"0A7F",
		X"0B50",
		X"0BF7",
		X"0CC8",
		X"0D6F",
		X"0E40",
		X"0EE7",
		X"0FB8",
		X"105F",
		X"1130",
		X"11D7",
		X"12A8",
		X"134F",
		X"1420",
		X"14C7",
		X"1598",
		X"163F",
		X"1710",
		X"17B7",
		X"1888",
		X"192F",
		X"1A00",
		X"1AA7",
		X"1B78",
		X"1C1F",
		X"1CF0",
		X"1D97",
		X"1E68",
		X"1F0F",
		X"1FE0",
		X"2087",
		X"2158",
		X"21FF",
		X"22D0",
		X"009F",
		X"0170",
		X"0217",
		X"02E8",
		X"038F",
		X"0460",
		X"0507",
		X"05D8",
		X"067F",
		X"0750",
		X"07F7",
		X"08C8",
		X"096F",
		X"0A40",
		X"0AE7",
		X"0BB8",
		X"0C5F",
		X"0D30",
		X"0DD7",
		X"0EA8",
		X"0F4F",
		X"1020",
		X"10C7",
		X"1198",
		X"123F",
		X"1310",
		X"13B7",
		X"1488",
		X"152F",
		X"1600",
		X"16A7",
		X"1778",
		X"181F",
		X"18F0",
		X"1997",
		X"1A68",
		X"1B0F",
		X"1BE0",
		X"1C87",
		X"1D58",
		X"1DFF",
		X"1ED0",
		X"1F77",
		X"2048",
		X"20EF",
		X"21C0",
		X"2267",
		X"0060",
		X"0107",
		X"01D8",
		X"027F",
		X"0350",
		X"03F7",
		X"04C8",
		X"056F",
		X"0640",
		X"06E7",
		X"07B8",
		X"085F",
		X"0930",
		X"09D7",
		X"0AA8",
		X"0B4F",
		X"0C20",
		X"0CC7",
		X"0D98",
		X"0E3F",
		X"0F10",
		X"0FB7",
		X"1088",
		X"112F",
		X"1200",
		X"12A7",
		X"1378",
		X"141F",
		X"14F0",
		X"1597",
		X"1668",
		X"170F",
		X"17E0",
		X"1887",
		X"1958",
		X"19FF",
		X"1AD0",
		X"1B77",
		X"1C48",
		X"1CEF",
		X"1DC0",
		X"1E67",
		X"1F38",
		X"1FDF",
		X"20B0",
		X"2157",
		X"2228",
		X"22CF",
		X"00C8",
		X"016F",
		X"0240",
		X"02E7",
		X"03B8",
		X"045F",
		X"0530",
		X"05D7",
		X"06A8",
		X"074F",
		X"0820",
		X"08C7",
		X"0998",
		X"0A3F",
		X"0B10",
		X"0BB7",
		X"0C88",
		X"0D2F",
		X"0E00",
		X"0EA7",
		X"0F78",
		X"101F",
		X"10F0",
		X"1197",
		X"1268",
		X"130F",
		X"13E0",
		X"1487",
		X"1558",
		X"15FF",
		X"16D0",
		X"1777",
		X"1848",
		X"18EF",
		X"19C0",
		X"1A67",
		X"1B38",
		X"1BDF",
		X"1CB0",
		X"1D57",
		X"1E28",
		X"1ECF",
		X"1FA0",
		X"2047",
		X"2118",
		X"21BF",
		X"2290",
		X"005F",
		X"0130",
		X"01D7",
		X"02A8",
		X"034F",
		X"0420",
		X"04C7",
		X"0598",
		X"063F",
		X"0710",
		X"07B7",
		X"0888",
		X"092F",
		X"0A00",
		X"0AA7",
		X"0B78",
		X"0C1F",
		X"0CF0",
		X"0D97",
		X"0E68",
		X"0F0F",
		X"0FE0",
		X"1087",
		X"1158",
		X"11FF",
		X"12D0",
		X"1377",
		X"1448",
		X"14EF",
		X"15C0",
		X"1667",
		X"1738",
		X"17DF",
		X"18B0",
		X"1957",
		X"1A28",
		X"1ACF",
		X"1BA0",
		X"1C47",
		X"1D18",
		X"1DBF",
		X"1E90",
		X"1F37",
		X"2008",
		X"20AF",
		X"2180",
		X"2227",
		X"0020",
		X"00C7",
		X"0198",
		X"023F",
		X"0310",
		X"03B7",
		X"0488",
		X"052F",
		X"0600",
		X"06A7",
		X"0778",
		X"081F",
		X"08F0",
		X"0997",
		X"0A68",
		X"0B0F",
		X"0BE0",
		X"0C87",
		X"0D58",
		X"0DFF",
		X"0ED0",
		X"0F77",
		X"1048",
		X"10EF",
		X"11C0",
		X"1267",
		X"1338",
		X"13DF",
		X"14B0",
		X"1557",
		X"1628",
		X"16CF",
		X"17A0",
		X"1847",
		X"1918",
		X"19BF",
		X"1A90",
		X"1B37",
		X"1C08",
		X"1CAF",
		X"1D80",
		X"1E27",
		X"1EF8",
		X"1F9F",
		X"2070",
		X"2117",
		X"21E8",
		X"228F",
		X"0088",
		X"012F",
		X"0200",
		X"02A7",
		X"0378",
		X"041F",
		X"04F0",
		X"0597",
		X"0668",
		X"070F",
		X"07E0",
		X"0887",
		X"0958",
		X"09FF",
		X"0AD0",
		X"0B77",
		X"0C48",
		X"0CEF",
		X"0DC0",
		X"0E67",
		X"0F38",
		X"0FDF",
		X"10B0",
		X"1157",
		X"1228",
		X"12CF",
		X"13A0",
		X"1447",
		X"1518",
		X"15BF",
		X"1690",
		X"1737",
		X"1808",
		X"18AF",
		X"1980",
		X"1A27",
		X"1AF8",
		X"1B9F",
		X"1C70",
		X"1D17",
		X"1DE8",
		X"1E8F",
		X"1F60",
		X"2007",
		X"20D8",
		X"217F",
		X"2250",
		X"001F",
		X"00F0",
		X"0197",
		X"0268",
		X"030F",
		X"03E0",
		X"0487",
		X"0558",
		X"05FF",
		X"06D0",
		X"0777",
		X"0848",
		X"08EF",
		X"09C0",
		X"0A67",
		X"0B38",
		X"0BDF",
		X"0CB0",
		X"0D57",
		X"0E28",
		X"0ECF",
		X"0FA0",
		X"1047",
		X"1118",
		X"11BF",
		X"1290",
		X"1337",
		X"1408",
		X"14AF",
		X"1580",
		X"1627",
		X"16F8",
		X"179F",
		X"1870",
		X"1917",
		X"19E8",
		X"1A8F",
		X"1B60",
		X"1C07",
		X"1CD8",
		X"1D7F",
		X"1E50",
		X"1EF7",
		X"1FC8",
		X"206F",
		X"2140",
		X"21E7",
		X"22B8",
		X"0087",
		X"0158",
		X"01FF",
		X"02D0",
		X"0377",
		X"0448",
		X"04EF",
		X"05C0",
		X"0667",
		X"0738",
		X"07DF",
		X"08B0",
		X"0957",
		X"0A28",
		X"0ACF",
		X"0BA0",
		X"0C47",
		X"0D18",
		X"0DBF",
		X"0E90",
		X"0F37",
		X"1008",
		X"10AF",
		X"1180",
		X"1227",
		X"12F8",
		X"139F",
		X"1470",
		X"1517",
		X"15E8",
		X"168F",
		X"1760",
		X"1807",
		X"18D8",
		X"197F",
		X"1A50",
		X"1AF7",
		X"1BC8",
		X"1C6F",
		X"1D40",
		X"1DE7",
		X"1EB8",
		X"1F5F",
		X"2030",
		X"20D7",
		X"21A8",
		X"224F",
		X"0048",
		X"00EF",
		X"01C0",
		X"0267",
		X"0338",
		X"03DF",
		X"04B0",
		X"0557",
		X"0628",
		X"06CF",
		X"07A0",
		X"0847",
		X"0918",
		X"09BF",
		X"0A90",
		X"0B37",
		X"0C08",
		X"0CAF",
		X"0D80",
		X"0E27",
		X"0EF8",
		X"0F9F",
		X"1070",
		X"1117",
		X"11E8",
		X"128F",
		X"1360",
		X"1407",
		X"14D8",
		X"157F",
		X"1650",
		X"16F7",
		X"17C8",
		X"186F",
		X"1940",
		X"19E7",
		X"1AB8",
		X"1B5F",
		X"1C30",
		X"1CD7",
		X"1DA8",
		X"1E4F",
		X"1F20",
		X"1FC7",
		X"2098",
		X"213F",
		X"2210",
		X"22B7",
		X"00B0",
		X"0157",
		X"0228",
		X"02CF",
		X"03A0",
		X"0447",
		X"0518",
		X"05BF",
		X"0690",
		X"0737",
		X"0808",
		X"08AF",
		X"0980",
		X"0A27",
		X"0AF8",
		X"0B9F",
		X"0C70",
		X"0D17",
		X"0DE8",
		X"0E8F",
		X"0F60",
		X"1007",
		X"10D8",
		X"117F",
		X"1250",
		X"12F7",
		X"13C8",
		X"146F",
		X"1540",
		X"15E7",
		X"16B8",
		X"175F",
		X"1830",
		X"18D7",
		X"19A8",
		X"1A4F",
		X"1B20",
		X"1BC7",
		X"1C98",
		X"1D3F",
		X"1E10",
		X"1EB7",
		X"1F88",
		X"202F",
		X"2100",
		X"21A7",
		X"2278",
		X"0047",
		X"0118",
		X"01BF",
		X"0290",
		X"0337",
		X"0408",
		X"04AF",
		X"0580",
		X"0627",
		X"06F8",
		X"079F",
		X"0870",
		X"0917",
		X"09E8",
		X"0A8F",
		X"0B60",
		X"0C07",
		X"0CD8",
		X"0D7F",
		X"0E50",
		X"0EF7",
		X"0FC8",
		X"106F",
		X"1140",
		X"11E7",
		X"12B8",
		X"135F",
		X"1430",
		X"14D7",
		X"15A8",
		X"164F",
		X"1720",
		X"17C7",
		X"1898",
		X"193F",
		X"1A10",
		X"1AB7",
		X"1B88",
		X"1C2F",
		X"1D00",
		X"1DA7",
		X"1E78",
		X"1F1F",
		X"1FF0",
		X"2097",
		X"2168",
		X"220F",
		X"0006",
		X"00AD",
		X"015E",
		X"0205",
		X"02B6",
		X"035D",
		X"040E",
		X"04B5",
		X"0566",
		X"060D",
		X"06BE",
		X"0765",
		X"0816",
		X"08BD",
		X"096E",
		X"0A15",
		X"0AC6",
		X"0B6D",
		X"0C1E",
		X"0CC5",
		X"0D76",
		X"0E1D",
		X"0ECE",
		X"0F75",
		X"1026",
		X"10CD",
		X"117E",
		X"1225",
		X"12D6",
		X"137D",
		X"142E",
		X"14D5",
		X"1586",
		X"162D",
		X"16DE",
		X"1785",
		X"1836",
		X"18DD",
		X"198E",
		X"1A35",
		X"1AE6",
		X"1B8D",
		X"1C3E",
		X"1CE5",
		X"1D96",
		X"1E3D",
		X"1EEE",
		X"1F95",
		X"2046",
		X"20ED",
		X"219E",
		X"2245",
		X"001E",
		X"00C5",
		X"0176",
		X"021D",
		X"02CE",
		X"0375",
		X"0426",
		X"04CD",
		X"057E",
		X"0625",
		X"06D6",
		X"077D",
		X"082E",
		X"08D5",
		X"0986",
		X"0A2D",
		X"0ADE",
		X"0B85",
		X"0C36",
		X"0CDD",
		X"0D8E",
		X"0E35",
		X"0EE6",
		X"0F8D",
		X"103E",
		X"10E5",
		X"1196",
		X"123D",
		X"12EE",
		X"1395",
		X"1446",
		X"14ED",
		X"159E",
		X"1645",
		X"16F6",
		X"179D",
		X"184E",
		X"18F5",
		X"19A6",
		X"1A4D",
		X"1AFE",
		X"1BA5",
		X"1C56",
		X"1CFD",
		X"1DAE",
		X"1E55",
		X"1F06",
		X"1FAD",
		X"205E",
		X"2105",
		X"21B6",
		X"225D",
		X"0036",
		X"00DD",
		X"018E",
		X"0235",
		X"02E6",
		X"038D",
		X"043E",
		X"04E5",
		X"0596",
		X"063D",
		X"06EE",
		X"0795",
		X"0846",
		X"08ED",
		X"099E",
		X"0A45",
		X"0AF6",
		X"0B9D",
		X"0C4E",
		X"0CF5",
		X"0DA6",
		X"0E4D",
		X"0EFE",
		X"0FA5",
		X"1056",
		X"10FD",
		X"11AE",
		X"1255",
		X"1306",
		X"13AD",
		X"145E",
		X"1505",
		X"15B6",
		X"165D",
		X"170E",
		X"17B5",
		X"1866",
		X"190D",
		X"19BE",
		X"1A65",
		X"1B16",
		X"1BBD",
		X"1C6E",
		X"1D15",
		X"1DC6",
		X"1E6D",
		X"1F1E",
		X"1FC5",
		X"2076",
		X"211D",
		X"21CE",
		X"2275",
		X"004E",
		X"00F5",
		X"01A6",
		X"024D",
		X"02FE",
		X"03A5",
		X"0456",
		X"04FD",
		X"05AE",
		X"0655",
		X"0706",
		X"07AD",
		X"085E",
		X"0905",
		X"09B6",
		X"0A5D",
		X"0B0E",
		X"0BB5",
		X"0C66",
		X"0D0D",
		X"0DBE",
		X"0E65",
		X"0F16",
		X"0FBD",
		X"106E",
		X"1115",
		X"11C6",
		X"126D",
		X"131E",
		X"13C5",
		X"1476",
		X"151D",
		X"15CE",
		X"1675",
		X"1726",
		X"17CD",
		X"187E",
		X"1925",
		X"19D6",
		X"1A7D",
		X"1B2E",
		X"1BD5",
		X"1C86",
		X"1D2D",
		X"1DDE",
		X"1E85",
		X"1F36",
		X"1FDD",
		X"208E",
		X"2135",
		X"21E6",
		X"228D",
		X"0066",
		X"010D",
		X"01BE",
		X"0265",
		X"0316",
		X"03BD",
		X"046E",
		X"0515",
		X"05C6",
		X"066D",
		X"071E",
		X"07C5",
		X"0876",
		X"091D",
		X"09CE",
		X"0A75",
		X"0B26",
		X"0BCD",
		X"0C7E",
		X"0D25",
		X"0DD6",
		X"0E7D",
		X"0F2E",
		X"0FD5",
		X"1086",
		X"112D",
		X"11DE",
		X"1285",
		X"1336",
		X"13DD",
		X"148E",
		X"1535",
		X"15E6",
		X"168D",
		X"173E",
		X"17E5",
		X"1896",
		X"193D",
		X"19EE",
		X"1A95",
		X"1B46",
		X"1BED",
		X"1C9E",
		X"1D45",
		X"1DF6",
		X"1E9D",
		X"1F4E",
		X"1FF5",
		X"20A6",
		X"214D",
		X"21FE",
		X"22A5",
		X"007E",
		X"0125",
		X"01D6",
		X"027D",
		X"032E",
		X"03D5",
		X"0486",
		X"052D",
		X"05DE",
		X"0685",
		X"0736",
		X"07DD",
		X"088E",
		X"0935",
		X"09E6",
		X"0A8D",
		X"0B3E",
		X"0BE5",
		X"0C96",
		X"0D3D",
		X"0DEE",
		X"0E95",
		X"0F46",
		X"0FED",
		X"109E",
		X"1145",
		X"11F6",
		X"129D",
		X"134E",
		X"13F5",
		X"14A6",
		X"154D",
		X"15FE",
		X"16A5",
		X"1756",
		X"17FD",
		X"18AE",
		X"1955",
		X"1A06",
		X"1AAD",
		X"1B5E",
		X"1C05",
		X"1CB6",
		X"1D5D",
		X"1E0E",
		X"1EB5",
		X"1F66",
		X"200D",
		X"20BE",
		X"2165",
		X"2216",
		X"22BD",
		X"0096",
		X"013D",
		X"01EE",
		X"0295",
		X"0346",
		X"03ED",
		X"049E",
		X"0545",
		X"05F6",
		X"069D",
		X"074E",
		X"07F5",
		X"08A6",
		X"094D",
		X"09FE",
		X"0AA5",
		X"0B56",
		X"0BFD",
		X"0CAE",
		X"0D55",
		X"0E06",
		X"0EAD",
		X"0F5E",
		X"1005",
		X"10B6",
		X"115D",
		X"120E",
		X"12B5",
		X"1366",
		X"140D",
		X"14BE",
		X"1565",
		X"1616",
		X"16BD",
		X"176E",
		X"1815",
		X"18C6",
		X"196D",
		X"1A1E",
		X"1AC5",
		X"1B76",
		X"1C1D",
		X"1CCE",
		X"1D75",
		X"1E26",
		X"1ECD",
		X"1F7E",
		X"2025",
		X"20D6",
		X"217D",
		X"222E",
		X"22D5",
		X"00AE",
		X"0155",
		X"0206",
		X"02AD",
		X"035E",
		X"0405",
		X"04B6",
		X"055D",
		X"060E",
		X"06B5",
		X"0766",
		X"080D",
		X"08BE",
		X"0965",
		X"0A16",
		X"0ABD",
		X"0B6E",
		X"0C15",
		X"0CC6",
		X"0D6D",
		X"0E1E",
		X"0EC5",
		X"0F76",
		X"101D",
		X"10CE",
		X"1175",
		X"1226",
		X"12CD",
		X"137E",
		X"1425",
		X"14D6",
		X"157D",
		X"162E",
		X"16D5",
		X"1786",
		X"182D",
		X"18DE",
		X"1985",
		X"1A36",
		X"1ADD",
		X"1B8E",
		X"1C35",
		X"1CE6",
		X"1D8D",
		X"1E3E",
		X"1EE5",
		X"1F96",
		X"203D",
		X"20EE",
		X"2195",
		X"2246",
		X"0015",
		X"00C6",
		X"016D",
		X"021E",
		X"02C5",
		X"0376",
		X"041D",
		X"04CE",
		X"0575",
		X"0626",
		X"06CD",
		X"077E",
		X"0825",
		X"08D6",
		X"097D",
		X"0A2E",
		X"0AD5",
		X"0B86",
		X"0C2D",
		X"0CDE",
		X"0D85",
		X"0E36",
		X"0EDD",
		X"0F8E",
		X"1035",
		X"10E6",
		X"118D",
		X"123E",
		X"12E5",
		X"1396",
		X"143D",
		X"14EE",
		X"1595",
		X"1646",
		X"16ED",
		X"179E",
		X"1845",
		X"18F6",
		X"199D",
		X"1A4E",
		X"1AF5",
		X"1BA6",
		X"1C4D",
		X"1CFE",
		X"1DA5",
		X"1E56",
		X"1EFD",
		X"1FAE",
		X"2055",
		X"2106",
		X"21AD",
		X"225E",
		X"002D",
		X"00DE",
		X"0185",
		X"0236",
		X"02DD",
		X"038E",
		X"0435",
		X"04E6",
		X"058D",
		X"063E",
		X"06E5",
		X"0796",
		X"083D",
		X"08EE",
		X"0995",
		X"0A46",
		X"0AED",
		X"0B9E",
		X"0C45",
		X"0CF6",
		X"0D9D",
		X"0E4E",
		X"0EF5",
		X"0FA6",
		X"104D",
		X"10FE",
		X"11A5",
		X"1256",
		X"12FD",
		X"13AE",
		X"1455",
		X"1506",
		X"15AD",
		X"165E",
		X"1705",
		X"17B6",
		X"185D",
		X"190E",
		X"19B5",
		X"1A66",
		X"1B0D",
		X"1BBE",
		X"1C65",
		X"1D16",
		X"1DBD",
		X"1E6E",
		X"1F15",
		X"1FC6",
		X"206D",
		X"211E",
		X"21C5",
		X"2276",
		X"0045",
		X"00F6",
		X"019D",
		X"024E",
		X"02F5",
		X"03A6",
		X"044D",
		X"04FE",
		X"05A5",
		X"0656",
		X"06FD",
		X"07AE",
		X"0855",
		X"0906",
		X"09AD",
		X"0A5E",
		X"0B05",
		X"0BB6",
		X"0C5D",
		X"0D0E",
		X"0DB5",
		X"0E66",
		X"0F0D",
		X"0FBE",
		X"1065",
		X"1116",
		X"11BD",
		X"126E",
		X"1315",
		X"13C6",
		X"146D",
		X"151E",
		X"15C5",
		X"1676",
		X"171D",
		X"17CE",
		X"1875",
		X"1926",
		X"19CD",
		X"1A7E",
		X"1B25",
		X"1BD6",
		X"1C7D",
		X"1D2E",
		X"1DD5",
		X"1E86",
		X"1F2D",
		X"1FDE",
		X"2085",
		X"2136",
		X"21DD",
		X"228E",
		X"005D",
		X"010E",
		X"01B5",
		X"0266",
		X"030D",
		X"03BE",
		X"0465",
		X"0516",
		X"05BD",
		X"066E",
		X"0715",
		X"07C6",
		X"086D",
		X"091E",
		X"09C5",
		X"0A76",
		X"0B1D",
		X"0BCE",
		X"0C75",
		X"0D26",
		X"0DCD",
		X"0E7E",
		X"0F25",
		X"0FD6",
		X"107D",
		X"112E",
		X"11D5",
		X"1286",
		X"132D",
		X"13DE",
		X"1485",
		X"1536",
		X"15DD",
		X"168E",
		X"1735",
		X"17E6",
		X"188D",
		X"193E",
		X"19E5",
		X"1A96",
		X"1B3D",
		X"1BEE",
		X"1C95",
		X"1D46",
		X"1DED",
		X"1E9E",
		X"1F45",
		X"1FF6",
		X"209D",
		X"214E",
		X"21F5",
		X"22A6",
		X"0075",
		X"0126",
		X"01CD",
		X"027E",
		X"0325",
		X"03D6",
		X"047D",
		X"052E",
		X"05D5",
		X"0686",
		X"072D",
		X"07DE",
		X"0885",
		X"0936",
		X"09DD",
		X"0A8E",
		X"0B35",
		X"0BE6",
		X"0C8D",
		X"0D3E",
		X"0DE5",
		X"0E96",
		X"0F3D",
		X"0FEE",
		X"1095",
		X"1146",
		X"11ED",
		X"129E",
		X"1345",
		X"13F6",
		X"149D",
		X"154E",
		X"15F5",
		X"16A6",
		X"174D",
		X"17FE",
		X"18A5",
		X"1956",
		X"19FD",
		X"1AAE",
		X"1B55",
		X"1C06",
		X"1CAD",
		X"1D5E",
		X"1E05",
		X"1EB6",
		X"1F5D",
		X"200E",
		X"20B5",
		X"2166",
		X"220D",
		X"22BE",
		X"008D",
		X"013E",
		X"01E5",
		X"0296",
		X"033D",
		X"03EE",
		X"0495",
		X"0546",
		X"05ED",
		X"069E",
		X"0745",
		X"07F6",
		X"089D",
		X"094E",
		X"09F5",
		X"0AA6",
		X"0B4D",
		X"0BFE",
		X"0CA5",
		X"0D56",
		X"0DFD",
		X"0EAE",
		X"0F55",
		X"1006",
		X"10AD",
		X"115E",
		X"1205",
		X"12B6",
		X"135D",
		X"140E",
		X"14B5",
		X"1566",
		X"160D",
		X"16BE",
		X"1765",
		X"1816",
		X"18BD",
		X"196E",
		X"1A15",
		X"1AC6",
		X"1B6D",
		X"1C1E",
		X"1CC5",
		X"1D76",
		X"1E1D",
		X"1ECE",
		X"1F75",
		X"2026",
		X"20CD",
		X"217E",
		X"2225",
		X"22D6",
		X"00A5",
		X"0156",
		X"01FD",
		X"02AE",
		X"0355",
		X"0406",
		X"04AD",
		X"055E",
		X"0605",
		X"06B6",
		X"075D",
		X"080E",
		X"08B5",
		X"0966",
		X"0A0D",
		X"0ABE",
		X"0B65",
		X"0C16",
		X"0CBD",
		X"0D6E",
		X"0E15",
		X"0EC6",
		X"0F6D",
		X"101E",
		X"10C5",
		X"1176",
		X"121D",
		X"12CE",
		X"1375",
		X"1426",
		X"14CD",
		X"157E",
		X"1625",
		X"16D6",
		X"177D",
		X"182E",
		X"18D5",
		X"1986",
		X"1A2D",
		X"1ADE",
		X"1B85",
		X"1C36",
		X"1CDD",
		X"1D8E",
		X"1E35",
		X"1EE6",
		X"1F8D",
		X"203E",
		X"20E5",
		X"2196",
		X"223D",
		X"0016",
		X"00BD",
		X"016E",
		X"0215",
		X"02C6",
		X"036D",
		X"041E",
		X"04C5",
		X"0576",
		X"061D",
		X"06CE",
		X"0775",
		X"0826",
		X"08CD",
		X"097E",
		X"0A25",
		X"0AD6",
		X"0B7D",
		X"0C2E",
		X"0CD5",
		X"0D86",
		X"0E2D",
		X"0EDE",
		X"0F85",
		X"1036",
		X"10DD",
		X"118E",
		X"1235",
		X"12E6",
		X"138D",
		X"143E",
		X"14E5",
		X"1596",
		X"163D",
		X"16EE",
		X"1795",
		X"1846",
		X"18ED",
		X"199E",
		X"1A45",
		X"1AF6",
		X"1B9D",
		X"1C4E",
		X"1CF5",
		X"1DA6",
		X"1E4D",
		X"1EFE",
		X"1FA5",
		X"2056",
		X"20FD",
		X"21AE",
		X"2255",
		X"002E",
		X"00D5",
		X"0186",
		X"022D",
		X"02DE",
		X"0385",
		X"0436",
		X"04DD",
		X"058E",
		X"0635",
		X"06E6",
		X"078D",
		X"083E",
		X"08E5",
		X"0996",
		X"0A3D",
		X"0AEE",
		X"0B95",
		X"0C46",
		X"0CED",
		X"0D9E",
		X"0E45",
		X"0EF6",
		X"0F9D",
		X"104E",
		X"10F5",
		X"11A6",
		X"124D",
		X"12FE",
		X"13A5",
		X"1456",
		X"14FD",
		X"15AE",
		X"1655",
		X"1706",
		X"17AD",
		X"185E",
		X"1905",
		X"19B6",
		X"1A5D",
		X"1B0E",
		X"1BB5",
		X"1C66",
		X"1D0D",
		X"1DBE",
		X"1E65",
		X"1F16",
		X"1FBD",
		X"206E",
		X"2115",
		X"21C6",
		X"226D",
		X"0046",
		X"00ED",
		X"019E",
		X"0245",
		X"02F6",
		X"039D",
		X"044E",
		X"04F5",
		X"05A6",
		X"064D",
		X"06FE",
		X"07A5",
		X"0856",
		X"08FD",
		X"09AE",
		X"0A55",
		X"0B06",
		X"0BAD",
		X"0C5E",
		X"0D05",
		X"0DB6",
		X"0E5D",
		X"0F0E",
		X"0FB5",
		X"1066",
		X"110D",
		X"11BE",
		X"1265",
		X"1316",
		X"13BD",
		X"146E",
		X"1515",
		X"15C6",
		X"166D",
		X"171E",
		X"17C5",
		X"1876",
		X"191D",
		X"19CE",
		X"1A75",
		X"1B26",
		X"1BCD",
		X"1C7E",
		X"1D25",
		X"1DD6",
		X"1E7D",
		X"1F2E",
		X"1FD5",
		X"2086",
		X"212D",
		X"21DE",
		X"2285",
		X"005E",
		X"0105",
		X"01B6",
		X"025D",
		X"030E",
		X"03B5",
		X"0466",
		X"050D",
		X"05BE",
		X"0665",
		X"0716",
		X"07BD",
		X"086E",
		X"0915",
		X"09C6",
		X"0A6D",
		X"0B1E",
		X"0BC5",
		X"0C76",
		X"0D1D",
		X"0DCE",
		X"0E75",
		X"0F26",
		X"0FCD",
		X"107E",
		X"1125",
		X"11D6",
		X"127D",
		X"132E",
		X"13D5",
		X"1486",
		X"152D",
		X"15DE",
		X"1685",
		X"1736",
		X"17DD",
		X"188E",
		X"1935",
		X"19E6",
		X"1A8D",
		X"1B3E",
		X"1BE5",
		X"1C96",
		X"1D3D",
		X"1DEE",
		X"1E95",
		X"1F46",
		X"1FED",
		X"209E",
		X"2145",
		X"21F6",
		X"229D",
		X"0076",
		X"011D",
		X"01CE",
		X"0275",
		X"0326",
		X"03CD",
		X"047E",
		X"0525",
		X"05D6",
		X"067D",
		X"072E",
		X"07D5",
		X"0886",
		X"092D",
		X"09DE",
		X"0A85",
		X"0B36",
		X"0BDD",
		X"0C8E",
		X"0D35",
		X"0DE6",
		X"0E8D",
		X"0F3E",
		X"0FE5",
		X"1096",
		X"113D",
		X"11EE",
		X"1295",
		X"1346",
		X"13ED",
		X"149E",
		X"1545",
		X"15F6",
		X"169D",
		X"174E",
		X"17F5",
		X"18A6",
		X"194D",
		X"19FE",
		X"1AA5",
		X"1B56",
		X"1BFD",
		X"1CAE",
		X"1D55",
		X"1E06",
		X"1EAD",
		X"1F5E",
		X"2005",
		X"20B6",
		X"215D",
		X"220E",
		X"22B5",
		X"008E",
		X"0135",
		X"01E6",
		X"028D",
		X"033E",
		X"03E5",
		X"0496",
		X"053D",
		X"05EE",
		X"0695",
		X"0746",
		X"07ED",
		X"089E",
		X"0945",
		X"09F6",
		X"0A9D",
		X"0B4E",
		X"0BF5",
		X"0CA6",
		X"0D4D",
		X"0DFE",
		X"0EA5",
		X"0F56",
		X"0FFD",
		X"10AE",
		X"1155",
		X"1206",
		X"12AD",
		X"135E",
		X"1405",
		X"14B6",
		X"155D",
		X"160E",
		X"16B5",
		X"1766",
		X"180D",
		X"18BE",
		X"1965",
		X"1A16",
		X"1ABD",
		X"1B6E",
		X"1C15",
		X"1CC6",
		X"1D6D",
		X"1E1E",
		X"1EC5",
		X"1F76",
		X"201D",
		X"20CE",
		X"2175",
		X"2226",
		X"22CD",
		X"00A6",
		X"014D",
		X"01FE",
		X"02A5",
		X"0356",
		X"03FD",
		X"04AE",
		X"0555",
		X"0606",
		X"06AD",
		X"075E",
		X"0805",
		X"08B6",
		X"095D",
		X"0A0E",
		X"0AB5",
		X"0B66",
		X"0C0D",
		X"0CBE",
		X"0D65",
		X"0E16",
		X"0EBD",
		X"0F6E",
		X"1015",
		X"10C6",
		X"116D",
		X"121E",
		X"12C5",
		X"1376",
		X"141D",
		X"14CE",
		X"1575",
		X"1626",
		X"16CD",
		X"177E",
		X"1825",
		X"18D6",
		X"197D",
		X"1A2E",
		X"1AD5",
		X"1B86",
		X"1C2D",
		X"1CDE",
		X"1D85",
		X"1E36",
		X"1EDD",
		X"1F8E",
		X"2035",
		X"20E6",
		X"218D",
		X"223E",
		X"000D",
		X"00BE",
		X"0165",
		X"0216",
		X"02BD",
		X"036E",
		X"0415",
		X"04C6",
		X"056D",
		X"061E",
		X"06C5",
		X"0776",
		X"081D",
		X"08CE",
		X"0975",
		X"0A26",
		X"0ACD",
		X"0B7E",
		X"0C25",
		X"0CD6",
		X"0D7D",
		X"0E2E",
		X"0ED5",
		X"0F86",
		X"102D",
		X"10DE",
		X"1185",
		X"1236",
		X"12DD",
		X"138E",
		X"1435",
		X"14E6",
		X"158D",
		X"163E",
		X"16E5",
		X"1796",
		X"183D",
		X"18EE",
		X"1995",
		X"1A46",
		X"1AED",
		X"1B9E",
		X"1C45",
		X"1CF6",
		X"1D9D",
		X"1E4E",
		X"1EF5",
		X"1FA6",
		X"204D",
		X"20FE",
		X"21A5",
		X"2256",
		X"0025",
		X"00D6",
		X"017D",
		X"022E",
		X"02D5",
		X"0386",
		X"042D",
		X"04DE",
		X"0585",
		X"0636",
		X"06DD",
		X"078E",
		X"0835",
		X"08E6",
		X"098D",
		X"0A3E",
		X"0AE5",
		X"0B96",
		X"0C3D",
		X"0CEE",
		X"0D95",
		X"0E46",
		X"0EED",
		X"0F9E",
		X"1045",
		X"10F6",
		X"119D",
		X"124E",
		X"12F5",
		X"13A6",
		X"144D",
		X"14FE",
		X"15A5",
		X"1656",
		X"16FD",
		X"17AE",
		X"1855",
		X"1906",
		X"19AD",
		X"1A5E",
		X"1B05",
		X"1BB6",
		X"1C5D",
		X"1D0E",
		X"1DB5",
		X"1E66",
		X"1F0D",
		X"1FBE",
		X"2065",
		X"2116",
		X"21BD",
		X"226E",
		X"003D",
		X"00EE",
		X"0195",
		X"0246",
		X"02ED",
		X"039E",
		X"0445",
		X"04F6",
		X"059D",
		X"064E",
		X"06F5",
		X"07A6",
		X"084D",
		X"08FE",
		X"09A5",
		X"0A56",
		X"0AFD",
		X"0BAE",
		X"0C55",
		X"0D06",
		X"0DAD",
		X"0E5E",
		X"0F05",
		X"0FB6",
		X"105D",
		X"110E",
		X"11B5",
		X"1266",
		X"130D",
		X"13BE",
		X"1465",
		X"1516",
		X"15BD",
		X"166E",
		X"1715",
		X"17C6",
		X"186D",
		X"191E",
		X"19C5",
		X"1A76",
		X"1B1D",
		X"1BCE",
		X"1C75",
		X"1D26",
		X"1DCD",
		X"1E7E",
		X"1F25",
		X"1FD6",
		X"207D",
		X"212E",
		X"21D5",
		X"2286",
		X"0055",
		X"0106",
		X"01AD",
		X"025E",
		X"0305",
		X"03B6",
		X"045D",
		X"050E",
		X"05B5",
		X"0666",
		X"070D",
		X"07BE",
		X"0865",
		X"0916",
		X"09BD",
		X"0A6E",
		X"0B15",
		X"0BC6",
		X"0C6D",
		X"0D1E",
		X"0DC5",
		X"0E76",
		X"0F1D",
		X"0FCE",
		X"1075",
		X"1126",
		X"11CD",
		X"127E",
		X"1325",
		X"13D6",
		X"147D",
		X"152E",
		X"15D5",
		X"1686",
		X"172D",
		X"17DE",
		X"1885",
		X"1936",
		X"19DD",
		X"1A8E",
		X"1B35",
		X"1BE6",
		X"1C8D",
		X"1D3E",
		X"1DE5",
		X"1E96",
		X"1F3D",
		X"1FEE",
		X"2095",
		X"2146",
		X"21ED",
		X"229E",
		X"006D",
		X"011E",
		X"01C5",
		X"0276",
		X"031D",
		X"03CE",
		X"0475",
		X"0526",
		X"05CD",
		X"067E",
		X"0725",
		X"07D6",
		X"087D",
		X"092E",
		X"09D5",
		X"0A86",
		X"0B2D",
		X"0BDE",
		X"0C85",
		X"0D36",
		X"0DDD",
		X"0E8E",
		X"0F35",
		X"0FE6",
		X"108D",
		X"113E",
		X"11E5",
		X"1296",
		X"133D",
		X"13EE",
		X"1495",
		X"1546",
		X"15ED",
		X"169E",
		X"1745",
		X"17F6",
		X"189D",
		X"194E",
		X"19F5",
		X"1AA6",
		X"1B4D",
		X"1BFE",
		X"1CA5",
		X"1D56",
		X"1DFD",
		X"1EAE",
		X"1F55",
		X"2006",
		X"20AD",
		X"215E",
		X"2205",
		X"22B6",
		X"0085",
		X"0136",
		X"01DD",
		X"028E",
		X"0335",
		X"03E6",
		X"048D",
		X"053E",
		X"05E5",
		X"0696",
		X"073D",
		X"07EE",
		X"0895",
		X"0946",
		X"09ED",
		X"0A9E",
		X"0B45",
		X"0BF6",
		X"0C9D",
		X"0D4E",
		X"0DF5",
		X"0EA6",
		X"0F4D",
		X"0FFE",
		X"10A5",
		X"1156",
		X"11FD",
		X"12AE",
		X"1355",
		X"1406",
		X"14AD",
		X"155E",
		X"1605",
		X"16B6",
		X"175D",
		X"180E",
		X"18B5",
		X"1966",
		X"1A0D",
		X"1ABE",
		X"1B65",
		X"1C16",
		X"1CBD",
		X"1D6E",
		X"1E15",
		X"1EC6",
		X"1F6D",
		X"201E",
		X"20C5",
		X"2176",
		X"221D",
		X"22CE",
		X"009D",
		X"014E",
		X"01F5",
		X"02A6",
		X"034D",
		X"03FE",
		X"04A5",
		X"0556",
		X"05FD",
		X"06AE",
		X"0755",
		X"0806",
		X"08AD",
		X"095E",
		X"0A05",
		X"0AB6",
		X"0B5D",
		X"0C0E",
		X"0CB5",
		X"0D66",
		X"0E0D",
		X"0EBE",
		X"0F65",
		X"1016",
		X"10BD",
		X"116E",
		X"1215",
		X"12C6",
		X"136D",
		X"141E",
		X"14C5",
		X"1576",
		X"161D",
		X"16CE",
		X"1775",
		X"1826",
		X"18CD",
		X"197E",
		X"1A25",
		X"1AD6",
		X"1B7D",
		X"1C2E",
		X"1CD5",
		X"1D86",
		X"1E2D",
		X"1EDE",
		X"1F85",
		X"2036",
		X"20DD",
		X"218E",
		X"2235",
		X"000E",
		X"00B5",
		X"0166",
		X"020D",
		X"02BE",
		X"0365",
		X"0416",
		X"04BD",
		X"056E",
		X"0615",
		X"06C6",
		X"076D",
		X"081E",
		X"08C5",
		X"0976",
		X"0A1D",
		X"0ACE",
		X"0B75",
		X"0C26",
		X"0CCD",
		X"0D7E",
		X"0E25",
		X"0ED6",
		X"0F7D",
		X"102E",
		X"10D5",
		X"1186",
		X"122D",
		X"12DE",
		X"1385",
		X"1436",
		X"14DD",
		X"158E",
		X"1635",
		X"16E6",
		X"178D",
		X"183E",
		X"18E5",
		X"1996",
		X"1A3D",
		X"1AEE",
		X"1B95",
		X"1C46",
		X"1CED",
		X"1D9E",
		X"1E45",
		X"1EF6",
		X"1F9D",
		X"204E",
		X"20F5",
		X"21A6",
		X"224D",
		X"0026",
		X"00CD",
		X"017E",
		X"0225",
		X"02D6",
		X"037D",
		X"042E",
		X"04D5",
		X"0586",
		X"062D",
		X"06DE",
		X"0785",
		X"0836",
		X"08DD",
		X"098E",
		X"0A35",
		X"0AE6",
		X"0B8D",
		X"0C3E",
		X"0CE5",
		X"0D96",
		X"0E3D",
		X"0EEE",
		X"0F95",
		X"1046",
		X"10ED",
		X"119E",
		X"1245",
		X"12F6",
		X"139D",
		X"144E",
		X"14F5",
		X"15A6",
		X"164D",
		X"16FE",
		X"17A5",
		X"1856",
		X"18FD",
		X"19AE",
		X"1A55",
		X"1B06",
		X"1BAD",
		X"1C5E",
		X"1D05",
		X"1DB6",
		X"1E5D",
		X"1F0E",
		X"1FB5",
		X"2066",
		X"210D",
		X"21BE",
		X"2265",
		X"003E",
		X"00E5",
		X"0196",
		X"023D",
		X"02EE",
		X"0395",
		X"0446",
		X"04ED",
		X"059E",
		X"0645",
		X"06F6",
		X"079D",
		X"084E",
		X"08F5",
		X"09A6",
		X"0A4D",
		X"0AFE",
		X"0BA5",
		X"0C56",
		X"0CFD",
		X"0DAE",
		X"0E55",
		X"0F06",
		X"0FAD",
		X"105E",
		X"1105",
		X"11B6",
		X"125D",
		X"130E",
		X"13B5",
		X"1466",
		X"150D",
		X"15BE",
		X"1665",
		X"1716",
		X"17BD",
		X"186E",
		X"1915",
		X"19C6",
		X"1A6D",
		X"1B1E",
		X"1BC5",
		X"1C76",
		X"1D1D",
		X"1DCE",
		X"1E75",
		X"1F26",
		X"1FCD",
		X"207E",
		X"2125",
		X"21D6",
		X"227D",
		X"0056",
		X"00FD",
		X"01AE",
		X"0255",
		X"0306",
		X"03AD",
		X"045E",
		X"0505",
		X"05B6",
		X"065D",
		X"070E",
		X"07B5",
		X"0866",
		X"090D",
		X"09BE",
		X"0A65",
		X"0B16",
		X"0BBD",
		X"0C6E",
		X"0D15",
		X"0DC6",
		X"0E6D",
		X"0F1E",
		X"0FC5",
		X"1076",
		X"111D",
		X"11CE",
		X"1275",
		X"1326",
		X"13CD",
		X"147E",
		X"1525",
		X"15D6",
		X"167D",
		X"172E",
		X"17D5",
		X"1886",
		X"192D",
		X"19DE",
		X"1A85",
		X"1B36",
		X"1BDD",
		X"1C8E",
		X"1D35",
		X"1DE6",
		X"1E8D",
		X"1F3E",
		X"1FE5",
		X"2096",
		X"213D",
		X"21EE",
		X"2295",
		X"006E",
		X"0115",
		X"01C6",
		X"026D",
		X"031E",
		X"03C5",
		X"0476",
		X"051D",
		X"05CE",
		X"0675",
		X"0726",
		X"07CD",
		X"087E",
		X"0925",
		X"09D6",
		X"0A7D",
		X"0B2E",
		X"0BD5",
		X"0C86",
		X"0D2D",
		X"0DDE",
		X"0E85",
		X"0F36",
		X"0FDD",
		X"108E",
		X"1135",
		X"11E6",
		X"128D",
		X"133E",
		X"13E5",
		X"1496",
		X"153D",
		X"15EE",
		X"1695",
		X"1746",
		X"17ED",
		X"189E",
		X"1945",
		X"19F6",
		X"1A9D",
		X"1B4E",
		X"1BF5",
		X"1CA6",
		X"1D4D",
		X"1DFE",
		X"1EA5",
		X"1F56",
		X"1FFD",
		X"20AE",
		X"2155",
		X"2206",
		X"22AD",
		X"0086",
		X"012D",
		X"01DE",
		X"0285",
		X"0336",
		X"03DD",
		X"048E",
		X"0535",
		X"05E6",
		X"068D",
		X"073E",
		X"07E5",
		X"0896",
		X"093D",
		X"09EE",
		X"0A95",
		X"0B46",
		X"0BED",
		X"0C9E",
		X"0D45",
		X"0DF6",
		X"0E9D",
		X"0F4E",
		X"0FF5",
		X"10A6",
		X"114D",
		X"11FE",
		X"12A5",
		X"1356",
		X"13FD",
		X"14AE",
		X"1555",
		X"1606",
		X"16AD",
		X"175E",
		X"1805",
		X"18B6",
		X"195D",
		X"1A0E",
		X"1AB5",
		X"1B66",
		X"1C0D",
		X"1CBE",
		X"1D65",
		X"1E16",
		X"1EBD",
		X"1F6E",
		X"2015",
		X"20C6",
		X"216D",
		X"221E",
		X"22C5",
		X"009E",
		X"0145",
		X"01F6",
		X"029D",
		X"034E",
		X"03F5",
		X"04A6",
		X"054D",
		X"05FE",
		X"06A5",
		X"0756",
		X"07FD",
		X"08AE",
		X"0955",
		X"0A06",
		X"0AAD",
		X"0B5E",
		X"0C05",
		X"0CB6",
		X"0D5D",
		X"0E0E",
		X"0EB5",
		X"0F66",
		X"100D",
		X"10BE",
		X"1165",
		X"1216",
		X"12BD",
		X"136E",
		X"1415",
		X"14C6",
		X"156D",
		X"161E",
		X"16C5",
		X"1776",
		X"181D",
		X"18CE",
		X"1975",
		X"1A26",
		X"1ACD",
		X"1B7E",
		X"1C25",
		X"1CD6",
		X"1D7D",
		X"1E2E",
		X"1ED5",
		X"1F86",
		X"202D",
		X"20DE",
		X"2185",
		X"2236",
		X"0005",
		X"00B6",
		X"015D",
		X"020E",
		X"02B5",
		X"0366",
		X"040D",
		X"04BE",
		X"0565",
		X"0616",
		X"06BD",
		X"076E",
		X"0815",
		X"08C6",
		X"096D",
		X"0A1E",
		X"0AC5",
		X"0B76",
		X"0C1D",
		X"0CCE",
		X"0D75",
		X"0E26",
		X"0ECD",
		X"0F7E",
		X"1025",
		X"10D6",
		X"117D",
		X"122E",
		X"12D5",
		X"1386",
		X"142D",
		X"14DE",
		X"1585",
		X"1636",
		X"16DD",
		X"178E",
		X"1835",
		X"18E6",
		X"198D",
		X"1A3E",
		X"1AE5",
		X"1B96",
		X"1C3D",
		X"1CEE",
		X"1D95",
		X"1E46",
		X"1EED",
		X"1F9E",
		X"2045",
		X"20F6",
		X"219D",
		X"224E",
		X"001D",
		X"00CE",
		X"0175",
		X"0226",
		X"02CD",
		X"037E",
		X"0425",
		X"04D6",
		X"057D",
		X"062E",
		X"06D5",
		X"0786",
		X"082D",
		X"08DE",
		X"0985",
		X"0A36",
		X"0ADD",
		X"0B8E",
		X"0C35",
		X"0CE6",
		X"0D8D",
		X"0E3E",
		X"0EE5",
		X"0F96",
		X"103D",
		X"10EE",
		X"1195",
		X"1246",
		X"12ED",
		X"139E",
		X"1445",
		X"14F6",
		X"159D",
		X"164E",
		X"16F5",
		X"17A6",
		X"184D",
		X"18FE",
		X"19A5",
		X"1A56",
		X"1AFD",
		X"1BAE",
		X"1C55",
		X"1D06",
		X"1DAD",
		X"1E5E",
		X"1F05",
		X"1FB6",
		X"205D",
		X"210E",
		X"21B5",
		X"2266",
		X"0035",
		X"00E6",
		X"018D",
		X"023E",
		X"02E5",
		X"0396",
		X"043D",
		X"04EE",
		X"0595",
		X"0646",
		X"06ED",
		X"079E",
		X"0845",
		X"08F6",
		X"099D",
		X"0A4E",
		X"0AF5",
		X"0BA6",
		X"0C4D",
		X"0CFE",
		X"0DA5",
		X"0E56",
		X"0EFD",
		X"0FAE",
		X"1055",
		X"1106",
		X"11AD",
		X"125E",
		X"1305",
		X"13B6",
		X"145D",
		X"150E",
		X"15B5",
		X"1666",
		X"170D",
		X"17BE",
		X"1865",
		X"1916",
		X"19BD",
		X"1A6E",
		X"1B15",
		X"1BC6",
		X"1C6D",
		X"1D1E",
		X"1DC5",
		X"1E76",
		X"1F1D",
		X"1FCE",
		X"2075",
		X"2126",
		X"21CD",
		X"227E",
		X"004D",
		X"00FE",
		X"01A5",
		X"0256",
		X"02FD",
		X"03AE",
		X"0455",
		X"0506",
		X"05AD",
		X"065E",
		X"0705",
		X"07B6",
		X"085D",
		X"090E",
		X"09B5",
		X"0A66",
		X"0B0D",
		X"0BBE",
		X"0C65",
		X"0D16",
		X"0DBD",
		X"0E6E",
		X"0F15",
		X"0FC6",
		X"106D",
		X"111E",
		X"11C5",
		X"1276",
		X"131D",
		X"13CE",
		X"1475",
		X"1526",
		X"15CD",
		X"167E",
		X"1725",
		X"17D6",
		X"187D",
		X"192E",
		X"19D5",
		X"1A86",
		X"1B2D",
		X"1BDE",
		X"1C85",
		X"1D36",
		X"1DDD",
		X"1E8E",
		X"1F35",
		X"1FE6",
		X"208D",
		X"213E",
		X"21E5",
		X"2296",
		X"0065",
		X"0116",
		X"01BD",
		X"026E",
		X"0315",
		X"03C6",
		X"046D",
		X"051E",
		X"05C5",
		X"0676",
		X"071D",
		X"07CE",
		X"0875",
		X"0926",
		X"09CD",
		X"0A7E",
		X"0B25",
		X"0BD6",
		X"0C7D",
		X"0D2E",
		X"0DD5",
		X"0E86",
		X"0F2D",
		X"0FDE",
		X"1085",
		X"1136",
		X"11DD",
		X"128E",
		X"1335",
		X"13E6",
		X"148D",
		X"153E",
		X"15E5",
		X"1696",
		X"173D",
		X"17EE",
		X"1895",
		X"1946",
		X"19ED",
		X"1A9E",
		X"1B45",
		X"1BF6",
		X"1C9D",
		X"1D4E",
		X"1DF5",
		X"1EA6",
		X"1F4D",
		X"1FFE",
		X"20A5",
		X"2156",
		X"21FD",
		X"22AE",
		X"007D",
		X"012E",
		X"01D5",
		X"0286",
		X"032D",
		X"03DE",
		X"0485",
		X"0536",
		X"05DD",
		X"068E",
		X"0735",
		X"07E6",
		X"088D",
		X"093E",
		X"09E5",
		X"0A96",
		X"0B3D",
		X"0BEE",
		X"0C95",
		X"0D46",
		X"0DED",
		X"0E9E",
		X"0F45",
		X"0FF6",
		X"109D",
		X"114E",
		X"11F5",
		X"12A6",
		X"134D",
		X"13FE",
		X"14A5",
		X"1556",
		X"15FD",
		X"16AE",
		X"1755",
		X"1806",
		X"18AD",
		X"195E",
		X"1A05",
		X"1AB6",
		X"1B5D",
		X"1C0E",
		X"1CB5",
		X"1D66",
		X"1E0D",
		X"1EBE",
		X"1F65",
		X"2016",
		X"20BD",
		X"216E",
		X"2215",
		X"22C6",
		X"0095",
		X"0146",
		X"01ED",
		X"029E",
		X"0345",
		X"03F6",
		X"049D",
		X"054E",
		X"05F5",
		X"06A6",
		X"074D",
		X"07FE",
		X"08A5",
		X"0956",
		X"09FD",
		X"0AAE",
		X"0B55",
		X"0C06",
		X"0CAD",
		X"0D5E",
		X"0E05",
		X"0EB6",
		X"0F5D",
		X"100E",
		X"10B5",
		X"1166",
		X"120D",
		X"12BE",
		X"1365",
		X"1416",
		X"14BD",
		X"156E",
		X"1615",
		X"16C6",
		X"176D",
		X"181E",
		X"18C5",
		X"1976",
		X"1A1D",
		X"1ACE",
		X"1B75",
		X"1C26",
		X"1CCD",
		X"1D7E",
		X"1E25",
		X"1ED6",
		X"1F7D",
		X"202E",
		X"20D5",
		X"2186",
		X"222D");


begin
process(clk)
    variable addr_mod : integer;
begin
	if (rstn='0')then
		address_out1<= (others=>'0');
		address_out2<= (others=>'0');
		elsif rising_edge(clk) then
			-- Step 1: 取模运算（地址范围 0~8919）
			addr_mod := to_integer(unsigned(address_in1)) mod 8920;

			-- Step 2: 读取 ROM
			address_out2 <= rom_reg(8919-addr_mod)-'1';
			address_out1 <= address_in1;
    end if;
end process;
    -- process(clk)
    -- begin
        -- if rising_edge(clk) then
            -- -- 根据输入的address_in1，读取rom_reg数组对应位置的值，并赋给address_in2
            -- -- address_in1应该是16位宽，表示从0到8919的地址范围
            -- address_out2 <= rom_reg(to_integer(unsigned(address_in1))); 
        -- end if;
    -- end process;
   -- architecture body
end architecture_Index_rom;
